module Butterfly_Exp8_Mant23(
  input wire clk,
  input wire [31:0] in0_r,
  input wire [31:0] in0_i,
  input wire [31:0] in1_r,
  input wire [31:0] in1_i,
  input wire [31:0] twd_r,
  input wire [31:0] twd_i,
  output wire [127:0] out
);
  // lint_off MULTIPLY
  function automatic [47:0] umul48b_24b_x_24b (input reg [23:0] lhs, input reg [23:0] rhs);
    begin
      umul48b_24b_x_24b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_in0_r;
  reg [31:0] p0_in0_i;
  reg [31:0] p0_in1_r;
  reg [31:0] p0_in1_i;
  reg [31:0] p0_twd_r;
  reg [31:0] p0_twd_i;
  always_ff @ (posedge clk) begin
    p0_in0_r <= in0_r;
    p0_in0_i <= in0_i;
    p0_in1_r <= in1_r;
    p0_in1_i <= in1_i;
    p0_twd_r <= twd_r;
    p0_twd_i <= twd_i;
  end

  // ===== Pipe stage 1:
  wire [22:0] p1_in1_r_fraction__10_comb;
  wire [7:0] p1_in1_r_bexp__9_comb;
  wire [22:0] p1_twd_r_fraction__10_comb;
  wire [7:0] p1_twd_r_bexp__9_comb;
  wire [22:0] p1_in1_i_fraction__10_comb;
  wire [7:0] p1_in1_i_bexp__9_comb;
  wire [22:0] p1_twd_i_fraction__10_comb;
  wire [7:0] p1_twd_i_bexp__9_comb;
  wire [23:0] p1_in1_r_fraction__11_comb;
  wire [23:0] p1_twd_r_fraction__11_comb;
  wire [23:0] p1_in1_i_fraction__11_comb;
  wire [23:0] p1_twd_i_fraction__11_comb;
  wire [8:0] p1_concat_7289_comb;
  wire [8:0] p1_concat_7290_comb;
  wire [23:0] p1_in1_r_fraction__12_comb;
  wire [23:0] p1_twd_r_fraction__12_comb;
  wire [8:0] p1_concat_7295_comb;
  wire [8:0] p1_concat_7296_comb;
  wire [23:0] p1_in1_i_fraction__12_comb;
  wire [23:0] p1_twd_i_fraction__12_comb;
  wire [8:0] p1_add_7302_comb;
  wire p1_eq_7303_comb;
  wire p1_eq_7304_comb;
  wire [47:0] p1_fraction__1_comb;
  wire [8:0] p1_add_7307_comb;
  wire p1_eq_7308_comb;
  wire p1_eq_7309_comb;
  wire [47:0] p1_fraction__8_comb;
  wire [8:0] p1_add_7312_comb;
  wire [47:0] p1_fraction__16_comb;
  wire [8:0] p1_add_7315_comb;
  wire [47:0] p1_fraction__24_comb;
  wire [9:0] p1_exp__1_comb;
  wire [47:0] p1_fraction__2_comb;
  wire [47:0] p1_sticky__1_comb;
  wire [9:0] p1_exp__4_comb;
  wire [47:0] p1_fraction__9_comb;
  wire [47:0] p1_sticky__2_comb;
  wire [9:0] p1_exp__8_comb;
  wire [47:0] p1_fraction__17_comb;
  wire [47:0] p1_sticky__4_comb;
  wire [9:0] p1_exp__12_comb;
  wire [47:0] p1_fraction__25_comb;
  wire [47:0] p1_sticky__6_comb;
  wire [9:0] p1_exp__2_comb;
  wire [47:0] p1_fraction__3_comb;
  wire [9:0] p1_exp__5_comb;
  wire [47:0] p1_fraction__10_comb;
  wire [9:0] p1_exp__9_comb;
  wire [47:0] p1_fraction__18_comb;
  wire [9:0] p1_exp__13_comb;
  wire [47:0] p1_fraction__26_comb;
  wire [9:0] p1_exp__3_comb;
  wire [9:0] p1_exp__6_comb;
  wire [9:0] p1_exp__10_comb;
  wire [9:0] p1_exp__14_comb;
  wire [47:0] p1_fraction__4_comb;
  wire [47:0] p1_sticky__5_comb;
  wire [47:0] p1_fraction__11_comb;
  wire [47:0] p1_sticky__3_comb;
  wire [47:0] p1_fraction__19_comb;
  wire [47:0] p1_sticky__7_comb;
  wire [47:0] p1_fraction__27_comb;
  wire [47:0] p1_sticky__8_comb;
  wire [47:0] p1_fraction__5_comb;
  wire [47:0] p1_fraction__12_comb;
  wire [47:0] p1_fraction__20_comb;
  wire [47:0] p1_fraction__28_comb;
  wire [22:0] p1_fraction__6_comb;
  wire [22:0] p1_fraction__13_comb;
  wire [22:0] p1_fraction__21_comb;
  wire [22:0] p1_fraction__29_comb;
  wire p1_greater_than_half_way__2_comb;
  wire [23:0] p1_fraction__7_comb;
  wire p1_greater_than_half_way__1_comb;
  wire [23:0] p1_fraction__14_comb;
  wire p1_greater_than_half_way__3_comb;
  wire [23:0] p1_fraction__22_comb;
  wire p1_greater_than_half_way__4_comb;
  wire [23:0] p1_fraction__30_comb;
  wire p1_do_round_up__2_comb;
  wire [23:0] p1_add_7470_comb;
  wire p1_do_round_up__1_comb;
  wire [23:0] p1_add_7472_comb;
  wire p1_do_round_up__3_comb;
  wire [23:0] p1_add_7474_comb;
  wire p1_do_round_up__4_comb;
  wire [23:0] p1_add_7476_comb;
  wire [23:0] p1_fraction__23_comb;
  wire [23:0] p1_fraction__15_comb;
  wire [23:0] p1_fraction__31_comb;
  wire [23:0] p1_fraction__32_comb;
  wire [9:0] p1_add_7486_comb;
  wire [9:0] p1_add_7488_comb;
  wire [9:0] p1_add_7490_comb;
  wire [9:0] p1_add_7492_comb;
  wire [9:0] p1_exp__11_comb;
  wire [9:0] p1_exp__7_comb;
  wire [9:0] p1_exp__15_comb;
  wire [9:0] p1_exp__16_comb;
  wire p1_sgt_7501_comb;
  wire p1_sgt_7502_comb;
  wire p1_sgt_7503_comb;
  wire p1_sgt_7504_comb;
  wire [8:0] p1_result_exp__1_comb;
  wire [7:0] p1_high_exp__3_comb;
  wire [7:0] p1_high_exp__4_comb;
  wire [8:0] p1_result_exp__2_comb;
  wire [7:0] p1_high_exp__6_comb;
  wire [7:0] p1_high_exp__1_comb;
  wire [8:0] p1_result_exp__6_comb;
  wire [8:0] p1_result_exp__9_comb;
  wire [8:0] p1_result_exp__4_comb;
  wire p1_eq_7522_comb;
  wire p1_eq_7524_comb;
  wire [8:0] p1_result_exp__3_comb;
  wire p1_eq_7527_comb;
  wire p1_eq_7529_comb;
  wire [8:0] p1_result_exp__7_comb;
  wire [8:0] p1_result_exp__10_comb;
  wire p1_and_7543_comb;
  wire p1_and_7544_comb;
  wire p1_and_7555_comb;
  wire p1_and_7556_comb;
  wire p1_has_0_arg__2_comb;
  wire p1_has_inf_arg__2_comb;
  wire p1_has_0_arg__1_comb;
  wire p1_has_inf_arg__1_comb;
  wire p1_has_0_arg__3_comb;
  wire p1_has_inf_arg__3_comb;
  wire p1_has_0_arg__4_comb;
  wire p1_has_inf_arg__4_comb;
  wire p1_nor_7593_comb;
  wire p1_and_7595_comb;
  wire p1_and_7596_comb;
  wire p1_nor_7598_comb;
  wire p1_and_7600_comb;
  wire p1_and_7601_comb;
  wire p1_nor_7603_comb;
  wire p1_nor_7606_comb;
  wire [22:0] p1_result_fraction__3_comb;
  wire p1_is_result_nan__2_comb;
  wire [22:0] p1_result_fraction__1_comb;
  wire p1_is_result_nan__1_comb;
  wire [22:0] p1_result_fraction__6_comb;
  wire p1_is_result_nan__3_comb;
  wire [22:0] p1_result_fraction__9_comb;
  wire p1_is_result_nan__4_comb;
  wire [22:0] p1_result_fraction__4_comb;
  wire [22:0] p1_nan_fraction__1_comb;
  wire [7:0] p1_high_exp__29_comb;
  wire [22:0] p1_result_fraction__2_comb;
  wire [22:0] p1_nan_fraction__5_comb;
  wire [7:0] p1_high_exp__28_comb;
  wire [22:0] p1_result_fraction__7_comb;
  wire [22:0] p1_nan_fraction__3_comb;
  wire [7:0] p1_high_exp__30_comb;
  wire [22:0] p1_result_fraction__10_comb;
  wire [22:0] p1_nan_fraction__4_comb;
  wire [7:0] p1_high_exp__31_comb;
  wire [22:0] p1_result_fraction__8_comb;
  wire [7:0] p1_result_exp__8_comb;
  wire [22:0] p1_result_fraction__5_comb;
  wire [7:0] p1_result_exp__5_comb;
  wire [22:0] p1_result_fraction__11_comb;
  wire [7:0] p1_result_exp__11_comb;
  wire [22:0] p1_result_fraction__12_comb;
  wire [7:0] p1_result_exp__12_comb;
  wire [5:0] p1_add_7688_comb;
  wire p1_ugt_7690_comb;
  wire [5:0] p1_add_7694_comb;
  wire [5:0] p1_add_7699_comb;
  wire p1_ugt_7701_comb;
  wire [5:0] p1_add_7705_comb;
  wire [27:0] p1_wide_x_comb;
  wire [7:0] p1_greater_exp_bexp_comb;
  wire [27:0] p1_wide_y_comb;
  wire [27:0] p1_wide_x__2_comb;
  wire [7:0] p1_greater_exp_bexp__1_comb;
  wire [27:0] p1_wide_y__2_comb;
  wire [27:0] p1_wide_x__1_comb;
  wire [7:0] p1_sub_7722_comb;
  wire [27:0] p1_wide_y__1_comb;
  wire [7:0] p1_sub_7724_comb;
  wire [27:0] p1_wide_x__3_comb;
  wire [7:0] p1_sub_7726_comb;
  wire [27:0] p1_wide_y__3_comb;
  wire [7:0] p1_sub_7728_comb;
  wire p1_in1_i_sign__2_comb;
  wire p1_twd_i_sign__2_comb;
  wire [27:0] p1_dropped_x_comb;
  wire [27:0] p1_dropped_y_comb;
  wire [27:0] p1_dropped_x__1_comb;
  wire [27:0] p1_dropped_y__1_comb;
  wire p1_result_sign__2_comb;
  wire p1_in1_r_sign__2_comb;
  wire p1_twd_r_sign__2_comb;
  wire p1_result_sign__3_comb;
  wire p1_result_sign__1_comb;
  wire [7:0] p1_shift_x_comb;
  wire p1_sticky_x_comb;
  wire [7:0] p1_shift_y_comb;
  wire p1_sticky_y_comb;
  wire p1_result_sign__6_comb;
  wire p1_result_sign__4_comb;
  wire [7:0] p1_shift_x__1_comb;
  wire p1_sticky_x__1_comb;
  wire [7:0] p1_shift_y__1_comb;
  wire p1_sticky_y__1_comb;
  wire p1_bd__1_sign_comb;
  wire p1_result_sign__5_comb;
  wire [27:0] p1_shifted_x_comb;
  wire [27:0] p1_shifted_y_comb;
  wire p1_result_sign__8_comb;
  wire p1_result_sign__7_comb;
  wire [27:0] p1_shifted_x__1_comb;
  wire [27:0] p1_shifted_y__1_comb;
  wire [7:0] p1_high_exp__32_comb;
  wire [7:0] p1_high_exp__33_comb;
  wire [7:0] p1_high_exp__34_comb;
  wire [7:0] p1_high_exp__35_comb;
  wire p1_greater_exp_sign_comb;
  wire [27:0] p1_addend_x_comb;
  wire [27:0] p1_addend_y_comb;
  wire p1_greater_exp_sign__1_comb;
  wire [27:0] p1_addend_x__2_comb;
  wire [27:0] p1_addend_y__2_comb;
  wire p1_eq_7818_comb;
  wire p1_eq_7819_comb;
  wire p1_eq_7820_comb;
  wire p1_eq_7821_comb;
  wire p1_eq_7822_comb;
  wire p1_eq_7823_comb;
  wire p1_eq_7824_comb;
  wire p1_eq_7825_comb;
  wire p1_and_7828_comb;
  wire p1_and_7829_comb;
  wire p1_and_7832_comb;
  wire p1_and_7833_comb;
  wire [27:0] p1_addend_x__1_comb;
  wire [27:0] p1_addend_y__1_comb;
  wire [27:0] p1_addend_x__3_comb;
  wire [27:0] p1_addend_y__3_comb;
  wire p1_has_pos_inf_comb;
  wire p1_has_neg_inf_comb;
  wire p1_has_pos_inf__1_comb;
  wire p1_has_neg_inf__1_comb;
  wire [28:0] p1_fraction__33_comb;
  wire [28:0] p1_fraction__34_comb;
  wire [27:0] p1_bit_slice_7802_comb;
  wire [27:0] p1_bit_slice_7803_comb;
  wire p1_bit_slice_7804_comb;
  wire p1_bit_slice_7805_comb;
  wire p1_ne_7808_comb;
  wire p1_ne_7809_comb;
  wire p1_nor_7854_comb;
  wire p1_nor_7858_comb;
  wire p1_is_result_nan__5_comb;
  wire p1_is_operand_inf_comb;
  wire p1_is_result_nan__6_comb;
  wire p1_is_operand_inf__1_comb;
  wire [22:0] p1_in0_r_fraction__6_comb;
  wire [7:0] p1_in0_r_bexp__6_comb;
  wire [22:0] p1_in0_i_fraction__6_comb;
  wire [7:0] p1_in0_i_bexp__6_comb;
  wire p1_fraction_is_zero_comb;
  wire p1_fraction_is_zero__1_comb;
  wire p1_not_7874_comb;
  wire p1_not_7875_comb;
  wire p1_in0_r_sign__2_comb;
  wire p1_in0_i_sign__2_comb;
  assign p1_in1_r_fraction__10_comb = p0_in1_r[22:0];
  assign p1_in1_r_bexp__9_comb = p0_in1_r[30:23];
  assign p1_twd_r_fraction__10_comb = p0_twd_r[22:0];
  assign p1_twd_r_bexp__9_comb = p0_twd_r[30:23];
  assign p1_in1_i_fraction__10_comb = p0_in1_i[22:0];
  assign p1_in1_i_bexp__9_comb = p0_in1_i[30:23];
  assign p1_twd_i_fraction__10_comb = p0_twd_i[22:0];
  assign p1_twd_i_bexp__9_comb = p0_twd_i[30:23];
  assign p1_in1_r_fraction__11_comb = {1'h0, p1_in1_r_fraction__10_comb} | 24'h80_0000;
  assign p1_twd_r_fraction__11_comb = {1'h0, p1_twd_r_fraction__10_comb} | 24'h80_0000;
  assign p1_in1_i_fraction__11_comb = {1'h0, p1_in1_i_fraction__10_comb} | 24'h80_0000;
  assign p1_twd_i_fraction__11_comb = {1'h0, p1_twd_i_fraction__10_comb} | 24'h80_0000;
  assign p1_concat_7289_comb = {1'h0, p1_in1_r_bexp__9_comb};
  assign p1_concat_7290_comb = {1'h0, p1_twd_r_bexp__9_comb};
  assign p1_in1_r_fraction__12_comb = p1_in1_r_fraction__11_comb & {24{p1_in1_r_bexp__9_comb != 8'h00}};
  assign p1_twd_r_fraction__12_comb = p1_twd_r_fraction__11_comb & {24{p1_twd_r_bexp__9_comb != 8'h00}};
  assign p1_concat_7295_comb = {1'h0, p1_in1_i_bexp__9_comb};
  assign p1_concat_7296_comb = {1'h0, p1_twd_i_bexp__9_comb};
  assign p1_in1_i_fraction__12_comb = p1_in1_i_fraction__11_comb & {24{p1_in1_i_bexp__9_comb != 8'h00}};
  assign p1_twd_i_fraction__12_comb = p1_twd_i_fraction__11_comb & {24{p1_twd_i_bexp__9_comb != 8'h00}};
  assign p1_add_7302_comb = p1_concat_7289_comb + p1_concat_7290_comb;
  assign p1_eq_7303_comb = p1_in1_r_bexp__9_comb == 8'h00;
  assign p1_eq_7304_comb = p1_twd_r_bexp__9_comb == 8'h00;
  assign p1_fraction__1_comb = umul48b_24b_x_24b(p1_in1_r_fraction__12_comb, p1_twd_r_fraction__12_comb);
  assign p1_add_7307_comb = p1_concat_7295_comb + p1_concat_7296_comb;
  assign p1_eq_7308_comb = p1_in1_i_bexp__9_comb == 8'h00;
  assign p1_eq_7309_comb = p1_twd_i_bexp__9_comb == 8'h00;
  assign p1_fraction__8_comb = umul48b_24b_x_24b(p1_in1_i_fraction__12_comb, p1_twd_i_fraction__12_comb);
  assign p1_add_7312_comb = p1_concat_7289_comb + p1_concat_7296_comb;
  assign p1_fraction__16_comb = umul48b_24b_x_24b(p1_in1_r_fraction__12_comb, p1_twd_i_fraction__12_comb);
  assign p1_add_7315_comb = p1_concat_7295_comb + p1_concat_7290_comb;
  assign p1_fraction__24_comb = umul48b_24b_x_24b(p1_in1_i_fraction__12_comb, p1_twd_r_fraction__12_comb);
  assign p1_exp__1_comb = {1'h0, p1_add_7302_comb} + 10'h381;
  assign p1_fraction__2_comb = p1_fraction__1_comb >> p1_fraction__1_comb[47];
  assign p1_sticky__1_comb = {47'h0000_0000_0000, p1_fraction__1_comb[0]};
  assign p1_exp__4_comb = {1'h0, p1_add_7307_comb} + 10'h381;
  assign p1_fraction__9_comb = p1_fraction__8_comb >> p1_fraction__8_comb[47];
  assign p1_sticky__2_comb = {47'h0000_0000_0000, p1_fraction__8_comb[0]};
  assign p1_exp__8_comb = {1'h0, p1_add_7312_comb} + 10'h381;
  assign p1_fraction__17_comb = p1_fraction__16_comb >> p1_fraction__16_comb[47];
  assign p1_sticky__4_comb = {47'h0000_0000_0000, p1_fraction__16_comb[0]};
  assign p1_exp__12_comb = {1'h0, p1_add_7315_comb} + 10'h381;
  assign p1_fraction__25_comb = p1_fraction__24_comb >> p1_fraction__24_comb[47];
  assign p1_sticky__6_comb = {47'h0000_0000_0000, p1_fraction__24_comb[0]};
  assign p1_exp__2_comb = p1_exp__1_comb & {10{~(p1_eq_7303_comb | p1_eq_7304_comb)}};
  assign p1_fraction__3_comb = p1_fraction__2_comb | p1_sticky__1_comb;
  assign p1_exp__5_comb = p1_exp__4_comb & {10{~(p1_eq_7308_comb | p1_eq_7309_comb)}};
  assign p1_fraction__10_comb = p1_fraction__9_comb | p1_sticky__2_comb;
  assign p1_exp__9_comb = p1_exp__8_comb & {10{~(p1_eq_7303_comb | p1_eq_7309_comb)}};
  assign p1_fraction__18_comb = p1_fraction__17_comb | p1_sticky__4_comb;
  assign p1_exp__13_comb = p1_exp__12_comb & {10{~(p1_eq_7308_comb | p1_eq_7304_comb)}};
  assign p1_fraction__26_comb = p1_fraction__25_comb | p1_sticky__6_comb;
  assign p1_exp__3_comb = p1_exp__2_comb + {9'h000, p1_fraction__1_comb[47]};
  assign p1_exp__6_comb = p1_exp__5_comb + {9'h000, p1_fraction__8_comb[47]};
  assign p1_exp__10_comb = p1_exp__9_comb + {9'h000, p1_fraction__16_comb[47]};
  assign p1_exp__14_comb = p1_exp__13_comb + {9'h000, p1_fraction__24_comb[47]};
  assign p1_fraction__4_comb = $signed(p1_exp__3_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__3_comb[47:1]} : p1_fraction__3_comb;
  assign p1_sticky__5_comb = {47'h0000_0000_0000, p1_fraction__3_comb[0]};
  assign p1_fraction__11_comb = $signed(p1_exp__6_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__10_comb[47:1]} : p1_fraction__10_comb;
  assign p1_sticky__3_comb = {47'h0000_0000_0000, p1_fraction__10_comb[0]};
  assign p1_fraction__19_comb = $signed(p1_exp__10_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__18_comb[47:1]} : p1_fraction__18_comb;
  assign p1_sticky__7_comb = {47'h0000_0000_0000, p1_fraction__18_comb[0]};
  assign p1_fraction__27_comb = $signed(p1_exp__14_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__26_comb[47:1]} : p1_fraction__26_comb;
  assign p1_sticky__8_comb = {47'h0000_0000_0000, p1_fraction__26_comb[0]};
  assign p1_fraction__5_comb = p1_fraction__4_comb | p1_sticky__5_comb;
  assign p1_fraction__12_comb = p1_fraction__11_comb | p1_sticky__3_comb;
  assign p1_fraction__20_comb = p1_fraction__19_comb | p1_sticky__7_comb;
  assign p1_fraction__28_comb = p1_fraction__27_comb | p1_sticky__8_comb;
  assign p1_fraction__6_comb = p1_fraction__5_comb[45:23];
  assign p1_fraction__13_comb = p1_fraction__12_comb[45:23];
  assign p1_fraction__21_comb = p1_fraction__20_comb[45:23];
  assign p1_fraction__29_comb = p1_fraction__28_comb[45:23];
  assign p1_greater_than_half_way__2_comb = p1_fraction__5_comb[22] & p1_fraction__5_comb[21:0] != 22'h00_0000;
  assign p1_fraction__7_comb = {1'h0, p1_fraction__6_comb};
  assign p1_greater_than_half_way__1_comb = p1_fraction__12_comb[22] & p1_fraction__12_comb[21:0] != 22'h00_0000;
  assign p1_fraction__14_comb = {1'h0, p1_fraction__13_comb};
  assign p1_greater_than_half_way__3_comb = p1_fraction__20_comb[22] & p1_fraction__20_comb[21:0] != 22'h00_0000;
  assign p1_fraction__22_comb = {1'h0, p1_fraction__21_comb};
  assign p1_greater_than_half_way__4_comb = p1_fraction__28_comb[22] & p1_fraction__28_comb[21:0] != 22'h00_0000;
  assign p1_fraction__30_comb = {1'h0, p1_fraction__29_comb};
  assign p1_do_round_up__2_comb = p1_greater_than_half_way__2_comb | p1_fraction__5_comb[22] & p1_fraction__5_comb[21:0] == 22'h00_0000 & p1_fraction__5_comb[23];
  assign p1_add_7470_comb = p1_fraction__7_comb + 24'h00_0001;
  assign p1_do_round_up__1_comb = p1_greater_than_half_way__1_comb | p1_fraction__12_comb[22] & p1_fraction__12_comb[21:0] == 22'h00_0000 & p1_fraction__12_comb[23];
  assign p1_add_7472_comb = p1_fraction__14_comb + 24'h00_0001;
  assign p1_do_round_up__3_comb = p1_greater_than_half_way__3_comb | p1_fraction__20_comb[22] & p1_fraction__20_comb[21:0] == 22'h00_0000 & p1_fraction__20_comb[23];
  assign p1_add_7474_comb = p1_fraction__22_comb + 24'h00_0001;
  assign p1_do_round_up__4_comb = p1_greater_than_half_way__4_comb | p1_fraction__28_comb[22] & p1_fraction__28_comb[21:0] == 22'h00_0000 & p1_fraction__28_comb[23];
  assign p1_add_7476_comb = p1_fraction__30_comb + 24'h00_0001;
  assign p1_fraction__23_comb = p1_do_round_up__2_comb ? p1_add_7470_comb : p1_fraction__7_comb;
  assign p1_fraction__15_comb = p1_do_round_up__1_comb ? p1_add_7472_comb : p1_fraction__14_comb;
  assign p1_fraction__31_comb = p1_do_round_up__3_comb ? p1_add_7474_comb : p1_fraction__22_comb;
  assign p1_fraction__32_comb = p1_do_round_up__4_comb ? p1_add_7476_comb : p1_fraction__30_comb;
  assign p1_add_7486_comb = p1_exp__3_comb + 10'h001;
  assign p1_add_7488_comb = p1_exp__6_comb + 10'h001;
  assign p1_add_7490_comb = p1_exp__10_comb + 10'h001;
  assign p1_add_7492_comb = p1_exp__14_comb + 10'h001;
  assign p1_exp__11_comb = p1_fraction__23_comb[23] ? p1_add_7486_comb : p1_exp__3_comb;
  assign p1_exp__7_comb = p1_fraction__15_comb[23] ? p1_add_7488_comb : p1_exp__6_comb;
  assign p1_exp__15_comb = p1_fraction__31_comb[23] ? p1_add_7490_comb : p1_exp__10_comb;
  assign p1_exp__16_comb = p1_fraction__32_comb[23] ? p1_add_7492_comb : p1_exp__14_comb;
  assign p1_sgt_7501_comb = $signed(p1_exp__11_comb) > $signed(10'h000);
  assign p1_sgt_7502_comb = $signed(p1_exp__7_comb) > $signed(10'h000);
  assign p1_sgt_7503_comb = $signed(p1_exp__15_comb) > $signed(10'h000);
  assign p1_sgt_7504_comb = $signed(p1_exp__16_comb) > $signed(10'h000);
  assign p1_result_exp__1_comb = p1_exp__11_comb[8:0];
  assign p1_high_exp__3_comb = 8'hff;
  assign p1_high_exp__4_comb = 8'hff;
  assign p1_result_exp__2_comb = p1_exp__7_comb[8:0];
  assign p1_high_exp__6_comb = 8'hff;
  assign p1_high_exp__1_comb = 8'hff;
  assign p1_result_exp__6_comb = p1_exp__15_comb[8:0];
  assign p1_result_exp__9_comb = p1_exp__16_comb[8:0];
  assign p1_result_exp__4_comb = p1_result_exp__1_comb & {9{p1_sgt_7501_comb}};
  assign p1_eq_7522_comb = p1_in1_r_bexp__9_comb == p1_high_exp__3_comb;
  assign p1_eq_7524_comb = p1_twd_r_bexp__9_comb == p1_high_exp__4_comb;
  assign p1_result_exp__3_comb = p1_result_exp__2_comb & {9{p1_sgt_7502_comb}};
  assign p1_eq_7527_comb = p1_in1_i_bexp__9_comb == p1_high_exp__6_comb;
  assign p1_eq_7529_comb = p1_twd_i_bexp__9_comb == p1_high_exp__1_comb;
  assign p1_result_exp__7_comb = p1_result_exp__6_comb & {9{p1_sgt_7503_comb}};
  assign p1_result_exp__10_comb = p1_result_exp__9_comb & {9{p1_sgt_7504_comb}};
  assign p1_and_7543_comb = p1_eq_7522_comb & p1_in1_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_7544_comb = p1_eq_7524_comb & p1_twd_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_7555_comb = p1_eq_7527_comb & p1_in1_i_fraction__10_comb == 23'h00_0000;
  assign p1_and_7556_comb = p1_eq_7529_comb & p1_twd_i_fraction__10_comb == 23'h00_0000;
  assign p1_has_0_arg__2_comb = p1_eq_7303_comb | p1_eq_7304_comb;
  assign p1_has_inf_arg__2_comb = p1_and_7543_comb | p1_and_7544_comb;
  assign p1_has_0_arg__1_comb = p1_eq_7308_comb | p1_eq_7309_comb;
  assign p1_has_inf_arg__1_comb = p1_and_7555_comb | p1_and_7556_comb;
  assign p1_has_0_arg__3_comb = p1_eq_7303_comb | p1_eq_7309_comb;
  assign p1_has_inf_arg__3_comb = p1_and_7543_comb | p1_and_7556_comb;
  assign p1_has_0_arg__4_comb = p1_eq_7308_comb | p1_eq_7304_comb;
  assign p1_has_inf_arg__4_comb = p1_and_7555_comb | p1_and_7544_comb;
  assign p1_nor_7593_comb = ~(p1_result_exp__4_comb[8] | p1_result_exp__4_comb[0] & p1_result_exp__4_comb[1] & p1_result_exp__4_comb[2] & p1_result_exp__4_comb[3] & p1_result_exp__4_comb[4] & p1_result_exp__4_comb[5] & p1_result_exp__4_comb[6] & p1_result_exp__4_comb[7]);
  assign p1_and_7595_comb = p1_eq_7522_comb & p1_in1_r_fraction__10_comb != 23'h00_0000;
  assign p1_and_7596_comb = p1_eq_7524_comb & p1_twd_r_fraction__10_comb != 23'h00_0000;
  assign p1_nor_7598_comb = ~(p1_result_exp__3_comb[8] | p1_result_exp__3_comb[0] & p1_result_exp__3_comb[1] & p1_result_exp__3_comb[2] & p1_result_exp__3_comb[3] & p1_result_exp__3_comb[4] & p1_result_exp__3_comb[5] & p1_result_exp__3_comb[6] & p1_result_exp__3_comb[7]);
  assign p1_and_7600_comb = p1_eq_7527_comb & p1_in1_i_fraction__10_comb != 23'h00_0000;
  assign p1_and_7601_comb = p1_eq_7529_comb & p1_twd_i_fraction__10_comb != 23'h00_0000;
  assign p1_nor_7603_comb = ~(p1_result_exp__7_comb[8] | p1_result_exp__7_comb[0] & p1_result_exp__7_comb[1] & p1_result_exp__7_comb[2] & p1_result_exp__7_comb[3] & p1_result_exp__7_comb[4] & p1_result_exp__7_comb[5] & p1_result_exp__7_comb[6] & p1_result_exp__7_comb[7]);
  assign p1_nor_7606_comb = ~(p1_result_exp__10_comb[8] | p1_result_exp__10_comb[0] & p1_result_exp__10_comb[1] & p1_result_exp__10_comb[2] & p1_result_exp__10_comb[3] & p1_result_exp__10_comb[4] & p1_result_exp__10_comb[5] & p1_result_exp__10_comb[6] & p1_result_exp__10_comb[7]);
  assign p1_result_fraction__3_comb = p1_fraction__23_comb[22:0];
  assign p1_is_result_nan__2_comb = p1_and_7595_comb | p1_and_7596_comb | p1_has_0_arg__2_comb & p1_has_inf_arg__2_comb;
  assign p1_result_fraction__1_comb = p1_fraction__15_comb[22:0];
  assign p1_is_result_nan__1_comb = p1_and_7600_comb | p1_and_7601_comb | p1_has_0_arg__1_comb & p1_has_inf_arg__1_comb;
  assign p1_result_fraction__6_comb = p1_fraction__31_comb[22:0];
  assign p1_is_result_nan__3_comb = p1_and_7595_comb | p1_and_7601_comb | p1_has_0_arg__3_comb & p1_has_inf_arg__3_comb;
  assign p1_result_fraction__9_comb = p1_fraction__32_comb[22:0];
  assign p1_is_result_nan__4_comb = p1_and_7600_comb | p1_and_7596_comb | p1_has_0_arg__4_comb & p1_has_inf_arg__4_comb;
  assign p1_result_fraction__4_comb = p1_result_fraction__3_comb & {23{p1_sgt_7501_comb}} & {23{p1_nor_7593_comb}} & {23{~(p1_and_7543_comb | p1_and_7544_comb)}};
  assign p1_nan_fraction__1_comb = 23'h40_0000;
  assign p1_high_exp__29_comb = 8'hff;
  assign p1_result_fraction__2_comb = p1_result_fraction__1_comb & {23{p1_sgt_7502_comb}} & {23{p1_nor_7598_comb}} & {23{~(p1_and_7555_comb | p1_and_7556_comb)}};
  assign p1_nan_fraction__5_comb = 23'h40_0000;
  assign p1_high_exp__28_comb = 8'hff;
  assign p1_result_fraction__7_comb = p1_result_fraction__6_comb & {23{p1_sgt_7503_comb}} & {23{p1_nor_7603_comb}} & {23{~(p1_and_7543_comb | p1_and_7556_comb)}};
  assign p1_nan_fraction__3_comb = 23'h40_0000;
  assign p1_high_exp__30_comb = 8'hff;
  assign p1_result_fraction__10_comb = p1_result_fraction__9_comb & {23{p1_sgt_7504_comb}} & {23{p1_nor_7606_comb}} & {23{~(p1_and_7555_comb | p1_and_7544_comb)}};
  assign p1_nan_fraction__4_comb = 23'h40_0000;
  assign p1_high_exp__31_comb = 8'hff;
  assign p1_result_fraction__8_comb = p1_is_result_nan__2_comb ? p1_nan_fraction__1_comb : p1_result_fraction__4_comb;
  assign p1_result_exp__8_comb = p1_is_result_nan__2_comb | p1_has_inf_arg__2_comb | ~p1_nor_7593_comb ? p1_high_exp__29_comb : p1_result_exp__4_comb[7:0];
  assign p1_result_fraction__5_comb = p1_is_result_nan__1_comb ? p1_nan_fraction__5_comb : p1_result_fraction__2_comb;
  assign p1_result_exp__5_comb = p1_is_result_nan__1_comb | p1_has_inf_arg__1_comb | ~p1_nor_7598_comb ? p1_high_exp__28_comb : p1_result_exp__3_comb[7:0];
  assign p1_result_fraction__11_comb = p1_is_result_nan__3_comb ? p1_nan_fraction__3_comb : p1_result_fraction__7_comb;
  assign p1_result_exp__11_comb = p1_is_result_nan__3_comb | p1_has_inf_arg__3_comb | ~p1_nor_7603_comb ? p1_high_exp__30_comb : p1_result_exp__7_comb[7:0];
  assign p1_result_fraction__12_comb = p1_is_result_nan__4_comb ? p1_nan_fraction__4_comb : p1_result_fraction__10_comb;
  assign p1_result_exp__12_comb = p1_is_result_nan__4_comb | p1_has_inf_arg__4_comb | ~p1_nor_7606_comb ? p1_high_exp__31_comb : p1_result_exp__10_comb[7:0];
  assign p1_add_7688_comb = p1_result_exp__8_comb[7:2] + 6'h07;
  assign p1_ugt_7690_comb = p1_result_exp__8_comb > p1_result_exp__5_comb;
  assign p1_add_7694_comb = p1_result_exp__5_comb[7:2] + 6'h07;
  assign p1_add_7699_comb = p1_result_exp__11_comb[7:2] + 6'h07;
  assign p1_ugt_7701_comb = p1_result_exp__11_comb > p1_result_exp__12_comb;
  assign p1_add_7705_comb = p1_result_exp__12_comb[7:2] + 6'h07;
  assign p1_wide_x_comb = {{2'h0, p1_result_fraction__8_comb} | 25'h080_0000, 3'h0};
  assign p1_greater_exp_bexp_comb = p1_ugt_7690_comb ? p1_result_exp__8_comb : p1_result_exp__5_comb;
  assign p1_wide_y_comb = {{2'h0, p1_result_fraction__5_comb} | 25'h080_0000, 3'h0};
  assign p1_wide_x__2_comb = {{2'h0, p1_result_fraction__11_comb} | 25'h080_0000, 3'h0};
  assign p1_greater_exp_bexp__1_comb = p1_ugt_7701_comb ? p1_result_exp__11_comb : p1_result_exp__12_comb;
  assign p1_wide_y__2_comb = {{2'h0, p1_result_fraction__12_comb} | 25'h080_0000, 3'h0};
  assign p1_wide_x__1_comb = p1_wide_x_comb & {28{p1_result_exp__8_comb != 8'h00}};
  assign p1_sub_7722_comb = {p1_add_7688_comb, p1_result_exp__8_comb[1:0]} - p1_greater_exp_bexp_comb;
  assign p1_wide_y__1_comb = p1_wide_y_comb & {28{p1_result_exp__5_comb != 8'h00}};
  assign p1_sub_7724_comb = {p1_add_7694_comb, p1_result_exp__5_comb[1:0]} - p1_greater_exp_bexp_comb;
  assign p1_wide_x__3_comb = p1_wide_x__2_comb & {28{p1_result_exp__11_comb != 8'h00}};
  assign p1_sub_7726_comb = {p1_add_7699_comb, p1_result_exp__11_comb[1:0]} - p1_greater_exp_bexp__1_comb;
  assign p1_wide_y__3_comb = p1_wide_y__2_comb & {28{p1_result_exp__12_comb != 8'h00}};
  assign p1_sub_7728_comb = {p1_add_7705_comb, p1_result_exp__12_comb[1:0]} - p1_greater_exp_bexp__1_comb;
  assign p1_in1_i_sign__2_comb = p0_in1_i[31:31];
  assign p1_twd_i_sign__2_comb = p0_twd_i[31:31];
  assign p1_dropped_x_comb = p1_sub_7722_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__1_comb << p1_sub_7722_comb;
  assign p1_dropped_y_comb = p1_sub_7724_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__1_comb << p1_sub_7724_comb;
  assign p1_dropped_x__1_comb = p1_sub_7726_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__3_comb << p1_sub_7726_comb;
  assign p1_dropped_y__1_comb = p1_sub_7728_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__3_comb << p1_sub_7728_comb;
  assign p1_result_sign__2_comb = p1_in1_i_sign__2_comb ^ p1_twd_i_sign__2_comb;
  assign p1_in1_r_sign__2_comb = p0_in1_r[31:31];
  assign p1_twd_r_sign__2_comb = p0_twd_r[31:31];
  assign p1_result_sign__3_comb = ~p1_is_result_nan__1_comb & p1_result_sign__2_comb;
  assign p1_result_sign__1_comb = p1_in1_r_sign__2_comb ^ p1_twd_r_sign__2_comb;
  assign p1_shift_x_comb = p1_greater_exp_bexp_comb - p1_result_exp__8_comb;
  assign p1_sticky_x_comb = p1_dropped_x_comb[27:3] != 25'h000_0000;
  assign p1_shift_y_comb = p1_greater_exp_bexp_comb - p1_result_exp__5_comb;
  assign p1_sticky_y_comb = p1_dropped_y_comb[27:3] != 25'h000_0000;
  assign p1_result_sign__6_comb = p1_in1_i_sign__2_comb ^ p1_twd_r_sign__2_comb;
  assign p1_result_sign__4_comb = p1_in1_r_sign__2_comb ^ p1_twd_i_sign__2_comb;
  assign p1_shift_x__1_comb = p1_greater_exp_bexp__1_comb - p1_result_exp__11_comb;
  assign p1_sticky_x__1_comb = p1_dropped_x__1_comb[27:3] != 25'h000_0000;
  assign p1_shift_y__1_comb = p1_greater_exp_bexp__1_comb - p1_result_exp__12_comb;
  assign p1_sticky_y__1_comb = p1_dropped_y__1_comb[27:3] != 25'h000_0000;
  assign p1_bd__1_sign_comb = ~p1_result_sign__3_comb;
  assign p1_result_sign__5_comb = ~p1_is_result_nan__2_comb & p1_result_sign__1_comb;
  assign p1_shifted_x_comb = p1_shift_x_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__1_comb >> p1_shift_x_comb;
  assign p1_shifted_y_comb = p1_shift_y_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__1_comb >> p1_shift_y_comb;
  assign p1_result_sign__8_comb = ~p1_is_result_nan__4_comb & p1_result_sign__6_comb;
  assign p1_result_sign__7_comb = ~p1_is_result_nan__3_comb & p1_result_sign__4_comb;
  assign p1_shifted_x__1_comb = p1_shift_x__1_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__3_comb >> p1_shift_x__1_comb;
  assign p1_shifted_y__1_comb = p1_shift_y__1_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__3_comb >> p1_shift_y__1_comb;
  assign p1_high_exp__32_comb = 8'hff;
  assign p1_high_exp__33_comb = 8'hff;
  assign p1_high_exp__34_comb = 8'hff;
  assign p1_high_exp__35_comb = 8'hff;
  assign p1_greater_exp_sign_comb = p1_ugt_7690_comb ? p1_result_sign__5_comb : p1_bd__1_sign_comb;
  assign p1_addend_x_comb = p1_shifted_x_comb | {27'h000_0000, p1_sticky_x_comb};
  assign p1_addend_y_comb = p1_shifted_y_comb | {27'h000_0000, p1_sticky_y_comb};
  assign p1_greater_exp_sign__1_comb = p1_ugt_7701_comb ? p1_result_sign__7_comb : p1_result_sign__8_comb;
  assign p1_addend_x__2_comb = p1_shifted_x__1_comb | {27'h000_0000, p1_sticky_x__1_comb};
  assign p1_addend_y__2_comb = p1_shifted_y__1_comb | {27'h000_0000, p1_sticky_y__1_comb};
  assign p1_eq_7818_comb = p1_result_exp__8_comb == p1_high_exp__32_comb;
  assign p1_eq_7819_comb = p1_result_fraction__8_comb == 23'h00_0000;
  assign p1_eq_7820_comb = p1_result_exp__5_comb == p1_high_exp__33_comb;
  assign p1_eq_7821_comb = p1_result_fraction__5_comb == 23'h00_0000;
  assign p1_eq_7822_comb = p1_result_exp__11_comb == p1_high_exp__34_comb;
  assign p1_eq_7823_comb = p1_result_fraction__11_comb == 23'h00_0000;
  assign p1_eq_7824_comb = p1_result_exp__12_comb == p1_high_exp__35_comb;
  assign p1_eq_7825_comb = p1_result_fraction__12_comb == 23'h00_0000;
  assign p1_and_7828_comb = p1_eq_7818_comb & p1_eq_7819_comb;
  assign p1_and_7829_comb = p1_eq_7820_comb & p1_eq_7821_comb;
  assign p1_and_7832_comb = p1_eq_7822_comb & p1_eq_7823_comb;
  assign p1_and_7833_comb = p1_eq_7824_comb & p1_eq_7825_comb;
  assign p1_addend_x__1_comb = p1_result_sign__5_comb ^ p1_greater_exp_sign_comb ? -p1_addend_x_comb : p1_addend_x_comb;
  assign p1_addend_y__1_comb = p1_bd__1_sign_comb ^ p1_greater_exp_sign_comb ? -p1_addend_y_comb : p1_addend_y_comb;
  assign p1_addend_x__3_comb = p1_result_sign__7_comb ^ p1_greater_exp_sign__1_comb ? -p1_addend_x__2_comb : p1_addend_x__2_comb;
  assign p1_addend_y__3_comb = p1_result_sign__8_comb ^ p1_greater_exp_sign__1_comb ? -p1_addend_y__2_comb : p1_addend_y__2_comb;
  assign p1_has_pos_inf_comb = ~(~(p1_eq_7818_comb & p1_eq_7819_comb) | p1_result_sign__5_comb) | ~(~(p1_eq_7820_comb & p1_eq_7821_comb) | p1_bd__1_sign_comb);
  assign p1_has_neg_inf_comb = p1_and_7828_comb & p1_result_sign__5_comb | p1_and_7829_comb & p1_bd__1_sign_comb;
  assign p1_has_pos_inf__1_comb = ~(~(p1_eq_7822_comb & p1_eq_7823_comb) | p1_result_sign__7_comb) | ~(~(p1_eq_7824_comb & p1_eq_7825_comb) | p1_result_sign__8_comb);
  assign p1_has_neg_inf__1_comb = p1_and_7832_comb & p1_result_sign__7_comb | p1_and_7833_comb & p1_result_sign__8_comb;
  assign p1_fraction__33_comb = {{1{p1_addend_x__1_comb[27]}}, p1_addend_x__1_comb} + {{1{p1_addend_y__1_comb[27]}}, p1_addend_y__1_comb};
  assign p1_fraction__34_comb = {{1{p1_addend_x__3_comb[27]}}, p1_addend_x__3_comb} + {{1{p1_addend_y__3_comb[27]}}, p1_addend_y__3_comb};
  assign p1_bit_slice_7802_comb = p1_fraction__33_comb[27:0];
  assign p1_bit_slice_7803_comb = p1_fraction__34_comb[27:0];
  assign p1_bit_slice_7804_comb = p1_fraction__33_comb[28];
  assign p1_bit_slice_7805_comb = p1_fraction__34_comb[28];
  assign p1_ne_7808_comb = p1_fraction__33_comb != 29'h0000_0000;
  assign p1_ne_7809_comb = p1_fraction__34_comb != 29'h0000_0000;
  assign p1_nor_7854_comb = ~(p1_and_7828_comb | p1_and_7829_comb);
  assign p1_nor_7858_comb = ~(p1_and_7832_comb | p1_and_7833_comb);
  assign p1_is_result_nan__5_comb = p1_eq_7818_comb & p1_result_fraction__8_comb != 23'h00_0000 | p1_eq_7820_comb & p1_result_fraction__5_comb != 23'h00_0000 | p1_has_pos_inf_comb & p1_has_neg_inf_comb;
  assign p1_is_operand_inf_comb = p1_and_7828_comb | p1_and_7829_comb;
  assign p1_is_result_nan__6_comb = p1_eq_7822_comb & p1_result_fraction__11_comb != 23'h00_0000 | p1_eq_7824_comb & p1_result_fraction__12_comb != 23'h00_0000 | p1_has_pos_inf__1_comb & p1_has_neg_inf__1_comb;
  assign p1_is_operand_inf__1_comb = p1_and_7832_comb | p1_and_7833_comb;
  assign p1_in0_r_fraction__6_comb = p0_in0_r[22:0];
  assign p1_in0_r_bexp__6_comb = p0_in0_r[30:23];
  assign p1_in0_i_fraction__6_comb = p0_in0_i[22:0];
  assign p1_in0_i_bexp__6_comb = p0_in0_i[30:23];
  assign p1_fraction_is_zero_comb = p1_fraction__33_comb == 29'h0000_0000;
  assign p1_fraction_is_zero__1_comb = p1_fraction__34_comb == 29'h0000_0000;
  assign p1_not_7874_comb = ~p1_has_pos_inf_comb;
  assign p1_not_7875_comb = ~p1_has_pos_inf__1_comb;
  assign p1_in0_r_sign__2_comb = p0_in0_r[31:31];
  assign p1_in0_i_sign__2_comb = p0_in0_i[31:31];

  // Registers for pipe stage 1:
  reg [7:0] p1_greater_exp_bexp;
  reg [7:0] p1_greater_exp_bexp__1;
  reg p1_greater_exp_sign;
  reg p1_greater_exp_sign__1;
  reg [27:0] p1_bit_slice_7802;
  reg [27:0] p1_bit_slice_7803;
  reg p1_bit_slice_7804;
  reg p1_bit_slice_7805;
  reg p1_ne_7808;
  reg p1_ne_7809;
  reg p1_nor_7854;
  reg p1_nor_7858;
  reg p1_is_result_nan__5;
  reg p1_is_operand_inf;
  reg p1_is_result_nan__6;
  reg p1_is_operand_inf__1;
  reg [22:0] p1_in0_r_fraction__6;
  reg [7:0] p1_in0_r_bexp__6;
  reg [22:0] p1_in0_i_fraction__6;
  reg [7:0] p1_in0_i_bexp__6;
  reg p1_fraction_is_zero;
  reg p1_fraction_is_zero__1;
  reg p1_not_7874;
  reg p1_not_7875;
  reg p1_in0_r_sign__2;
  reg p1_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p1_greater_exp_bexp <= p1_greater_exp_bexp_comb;
    p1_greater_exp_bexp__1 <= p1_greater_exp_bexp__1_comb;
    p1_greater_exp_sign <= p1_greater_exp_sign_comb;
    p1_greater_exp_sign__1 <= p1_greater_exp_sign__1_comb;
    p1_bit_slice_7802 <= p1_bit_slice_7802_comb;
    p1_bit_slice_7803 <= p1_bit_slice_7803_comb;
    p1_bit_slice_7804 <= p1_bit_slice_7804_comb;
    p1_bit_slice_7805 <= p1_bit_slice_7805_comb;
    p1_ne_7808 <= p1_ne_7808_comb;
    p1_ne_7809 <= p1_ne_7809_comb;
    p1_nor_7854 <= p1_nor_7854_comb;
    p1_nor_7858 <= p1_nor_7858_comb;
    p1_is_result_nan__5 <= p1_is_result_nan__5_comb;
    p1_is_operand_inf <= p1_is_operand_inf_comb;
    p1_is_result_nan__6 <= p1_is_result_nan__6_comb;
    p1_is_operand_inf__1 <= p1_is_operand_inf__1_comb;
    p1_in0_r_fraction__6 <= p1_in0_r_fraction__6_comb;
    p1_in0_r_bexp__6 <= p1_in0_r_bexp__6_comb;
    p1_in0_i_fraction__6 <= p1_in0_i_fraction__6_comb;
    p1_in0_i_bexp__6 <= p1_in0_i_bexp__6_comb;
    p1_fraction_is_zero <= p1_fraction_is_zero_comb;
    p1_fraction_is_zero__1 <= p1_fraction_is_zero__1_comb;
    p1_not_7874 <= p1_not_7874_comb;
    p1_not_7875 <= p1_not_7875_comb;
    p1_in0_r_sign__2 <= p1_in0_r_sign__2_comb;
    p1_in0_i_sign__2 <= p1_in0_i_sign__2_comb;
  end

  // ===== Pipe stage 2:
  wire [27:0] p2_abs_fraction_comb;
  wire [27:0] p2_abs_fraction__1_comb;
  wire [27:0] p2_reverse_7937_comb;
  wire [27:0] p2_reverse_7938_comb;
  wire [28:0] p2_one_hot_7939_comb;
  wire [28:0] p2_one_hot_7940_comb;
  wire [4:0] p2_encode_7941_comb;
  wire [4:0] p2_encode_7942_comb;
  wire p2_carry_bit_comb;
  wire p2_cancel_comb;
  wire p2_carry_bit__1_comb;
  wire p2_cancel__1_comb;
  wire [27:0] p2_leading_zeroes_comb;
  wire [27:0] p2_leading_zeroes__1_comb;
  wire p2_and_7969_comb;
  wire p2_and_7970_comb;
  wire p2_and_7971_comb;
  wire [26:0] p2_carry_fraction_comb;
  wire [27:0] p2_add_7975_comb;
  wire p2_and_7976_comb;
  wire p2_and_7977_comb;
  wire p2_and_7978_comb;
  wire [26:0] p2_carry_fraction__2_comb;
  wire [27:0] p2_add_7982_comb;
  wire [2:0] p2_concat_7983_comb;
  wire [26:0] p2_carry_fraction__1_comb;
  wire [26:0] p2_cancel_fraction_comb;
  wire [2:0] p2_concat_7986_comb;
  wire [26:0] p2_carry_fraction__3_comb;
  wire [26:0] p2_cancel_fraction__1_comb;
  wire [26:0] p2_shifted_fraction_comb;
  wire [26:0] p2_shifted_fraction__1_comb;
  wire [2:0] p2_normal_chunk_comb;
  wire [1:0] p2_half_way_chunk_comb;
  wire [2:0] p2_normal_chunk__1_comb;
  wire [1:0] p2_half_way_chunk__1_comb;
  wire [24:0] p2_add_8010_comb;
  wire [24:0] p2_add_8014_comb;
  wire p2_do_round_up__5_comb;
  wire p2_do_round_up__6_comb;
  wire [27:0] p2_rounded_fraction_comb;
  wire [27:0] p2_rounded_fraction__1_comb;
  wire p2_rounding_carry_comb;
  wire p2_rounding_carry__1_comb;
  wire [8:0] p2_add_8034_comb;
  wire [8:0] p2_add_8036_comb;
  wire [9:0] p2_add_8043_comb;
  wire [9:0] p2_add_8045_comb;
  wire [9:0] p2_wide_exponent_comb;
  wire [9:0] p2_wide_exponent__3_comb;
  wire [9:0] p2_wide_exponent__1_comb;
  wire [9:0] p2_wide_exponent__4_comb;
  wire [8:0] p2_wide_exponent__2_comb;
  wire [8:0] p2_wide_exponent__5_comb;
  wire [2:0] p2_add_8089_comb;
  wire [2:0] p2_add_8092_comb;
  wire [27:0] p2_shrl_8095_comb;
  wire p2_nor_8097_comb;
  wire [27:0] p2_shrl_8098_comb;
  wire p2_nor_8100_comb;
  wire [22:0] p2_result_fraction__13_comb;
  wire [22:0] p2_result_fraction__15_comb;
  wire [22:0] p2_result_fraction__14_comb;
  wire [22:0] p2_nan_fraction__14_comb;
  wire [7:0] p2_high_exp__36_comb;
  wire [22:0] p2_result_fraction__16_comb;
  wire [22:0] p2_nan_fraction__15_comb;
  wire [7:0] p2_high_exp__37_comb;
  wire [22:0] p2_result_fraction__17_comb;
  wire [7:0] p2_result_exponent__2_comb;
  wire [22:0] p2_result_fraction__18_comb;
  wire [7:0] p2_result_exponent__1_comb;
  wire [5:0] p2_add_8152_comb;
  wire p2_ugt_8154_comb;
  wire [5:0] p2_add_8163_comb;
  wire p2_ugt_8165_comb;
  wire p2_result_sign__9_comb;
  wire p2_result_sign__11_comb;
  wire [5:0] p2_add_8158_comb;
  wire [5:0] p2_add_8169_comb;
  wire [27:0] p2_wide_x__4_comb;
  wire [7:0] p2_greater_exp_bexp__2_comb;
  wire [27:0] p2_wide_x__6_comb;
  wire [7:0] p2_greater_exp_bexp__3_comb;
  wire [7:0] p2_high_exp__39_comb;
  wire p2_result_sign__10_comb;
  wire [7:0] p2_high_exp__41_comb;
  wire p2_result_sign__12_comb;
  wire [27:0] p2_wide_y__4_comb;
  wire [27:0] p2_wide_y__6_comb;
  wire [27:0] p2_wide_x__5_comb;
  wire [7:0] p2_sub_8190_comb;
  wire [27:0] p2_wide_x__7_comb;
  wire [7:0] p2_sub_8194_comb;
  wire [7:0] p2_high_exp__46_comb;
  wire p2_eq_8251_comb;
  wire p2_eq_8252_comb;
  wire [7:0] p2_high_exp__38_comb;
  wire p2_result_sign__13_comb;
  wire [7:0] p2_high_exp__47_comb;
  wire p2_eq_8257_comb;
  wire p2_eq_8258_comb;
  wire [7:0] p2_high_exp__40_comb;
  wire p2_result_sign__14_comb;
  wire [27:0] p2_wide_y__5_comb;
  wire [7:0] p2_sub_8192_comb;
  wire [27:0] p2_wide_y__7_comb;
  wire [7:0] p2_sub_8196_comb;
  wire [27:0] p2_dropped_x__2_comb;
  wire [27:0] p2_dropped_x__3_comb;
  wire p2_ne_8262_comb;
  wire p2_nand_8263_comb;
  wire p2_eq_8264_comb;
  wire p2_eq_8265_comb;
  wire p2_re__1_sign_comb;
  wire p2_ne_8267_comb;
  wire p2_nand_8268_comb;
  wire p2_eq_8269_comb;
  wire p2_eq_8270_comb;
  wire p2_im__1_sign_comb;
  wire [27:0] p2_dropped_y__2_comb;
  wire [27:0] p2_dropped_y__3_comb;
  wire p2_nor_8272_comb;
  wire p2_nor_8273_comb;
  wire p2_and_8274_comb;
  wire p2_nor_8275_comb;
  wire p2_nor_8277_comb;
  wire p2_nor_8278_comb;
  wire p2_and_8279_comb;
  wire p2_nor_8280_comb;
  wire [7:0] p2_shift_x__2_comb;
  wire p2_sticky_x__2_comb;
  wire [7:0] p2_shift_x__3_comb;
  wire p2_sticky_x__3_comb;
  wire p2_has_pos_inf__2_comb;
  wire p2_has_neg_inf__2_comb;
  wire p2_has_pos_inf__3_comb;
  wire p2_has_neg_inf__3_comb;
  wire p2_has_pos_inf__4_comb;
  wire p2_has_neg_inf__4_comb;
  wire p2_has_pos_inf__5_comb;
  wire p2_has_neg_inf__5_comb;
  wire [7:0] p2_shift_y__2_comb;
  wire p2_sticky_y__2_comb;
  wire [7:0] p2_shift_y__3_comb;
  wire p2_sticky_y__3_comb;
  wire [27:0] p2_shifted_x__2_comb;
  wire [27:0] p2_shifted_x__3_comb;
  wire p2_and_8284_comb;
  wire p2_and_8285_comb;
  wire p2_and_8289_comb;
  wire p2_and_8290_comb;
  wire p2_and_8295_comb;
  wire p2_and_8296_comb;
  wire p2_and_8299_comb;
  wire p2_and_8300_comb;
  wire [27:0] p2_shifted_y__2_comb;
  wire [27:0] p2_concat_8236_comb;
  wire [27:0] p2_shifted_y__3_comb;
  wire [27:0] p2_concat_8240_comb;
  wire [27:0] p2_addend_x__4_comb;
  wire [27:0] p2_addend_x__6_comb;
  wire p2_nor_8298_comb;
  wire p2_nor_8302_comb;
  wire p2_is_result_nan__7_comb;
  wire p2_is_operand_inf__2_comb;
  wire p2_not_8307_comb;
  wire p2_is_result_nan__8_comb;
  wire p2_is_operand_inf__3_comb;
  wire p2_not_8310_comb;
  wire p2_is_result_nan__9_comb;
  wire p2_not_8312_comb;
  wire p2_is_result_nan__10_comb;
  wire p2_not_8314_comb;
  assign p2_abs_fraction_comb = p1_bit_slice_7804 ? -p1_bit_slice_7802 : p1_bit_slice_7802;
  assign p2_abs_fraction__1_comb = p1_bit_slice_7805 ? -p1_bit_slice_7803 : p1_bit_slice_7803;
  assign p2_reverse_7937_comb = {p2_abs_fraction_comb[0], p2_abs_fraction_comb[1], p2_abs_fraction_comb[2], p2_abs_fraction_comb[3], p2_abs_fraction_comb[4], p2_abs_fraction_comb[5], p2_abs_fraction_comb[6], p2_abs_fraction_comb[7], p2_abs_fraction_comb[8], p2_abs_fraction_comb[9], p2_abs_fraction_comb[10], p2_abs_fraction_comb[11], p2_abs_fraction_comb[12], p2_abs_fraction_comb[13], p2_abs_fraction_comb[14], p2_abs_fraction_comb[15], p2_abs_fraction_comb[16], p2_abs_fraction_comb[17], p2_abs_fraction_comb[18], p2_abs_fraction_comb[19], p2_abs_fraction_comb[20], p2_abs_fraction_comb[21], p2_abs_fraction_comb[22], p2_abs_fraction_comb[23], p2_abs_fraction_comb[24], p2_abs_fraction_comb[25], p2_abs_fraction_comb[26], p2_abs_fraction_comb[27]};
  assign p2_reverse_7938_comb = {p2_abs_fraction__1_comb[0], p2_abs_fraction__1_comb[1], p2_abs_fraction__1_comb[2], p2_abs_fraction__1_comb[3], p2_abs_fraction__1_comb[4], p2_abs_fraction__1_comb[5], p2_abs_fraction__1_comb[6], p2_abs_fraction__1_comb[7], p2_abs_fraction__1_comb[8], p2_abs_fraction__1_comb[9], p2_abs_fraction__1_comb[10], p2_abs_fraction__1_comb[11], p2_abs_fraction__1_comb[12], p2_abs_fraction__1_comb[13], p2_abs_fraction__1_comb[14], p2_abs_fraction__1_comb[15], p2_abs_fraction__1_comb[16], p2_abs_fraction__1_comb[17], p2_abs_fraction__1_comb[18], p2_abs_fraction__1_comb[19], p2_abs_fraction__1_comb[20], p2_abs_fraction__1_comb[21], p2_abs_fraction__1_comb[22], p2_abs_fraction__1_comb[23], p2_abs_fraction__1_comb[24], p2_abs_fraction__1_comb[25], p2_abs_fraction__1_comb[26], p2_abs_fraction__1_comb[27]};
  assign p2_one_hot_7939_comb = {p2_reverse_7937_comb[27:0] == 28'h000_0000, p2_reverse_7937_comb[27] && p2_reverse_7937_comb[26:0] == 27'h000_0000, p2_reverse_7937_comb[26] && p2_reverse_7937_comb[25:0] == 26'h000_0000, p2_reverse_7937_comb[25] && p2_reverse_7937_comb[24:0] == 25'h000_0000, p2_reverse_7937_comb[24] && p2_reverse_7937_comb[23:0] == 24'h00_0000, p2_reverse_7937_comb[23] && p2_reverse_7937_comb[22:0] == 23'h00_0000, p2_reverse_7937_comb[22] && p2_reverse_7937_comb[21:0] == 22'h00_0000, p2_reverse_7937_comb[21] && p2_reverse_7937_comb[20:0] == 21'h00_0000, p2_reverse_7937_comb[20] && p2_reverse_7937_comb[19:0] == 20'h0_0000, p2_reverse_7937_comb[19] && p2_reverse_7937_comb[18:0] == 19'h0_0000, p2_reverse_7937_comb[18] && p2_reverse_7937_comb[17:0] == 18'h0_0000, p2_reverse_7937_comb[17] && p2_reverse_7937_comb[16:0] == 17'h0_0000, p2_reverse_7937_comb[16] && p2_reverse_7937_comb[15:0] == 16'h0000, p2_reverse_7937_comb[15] && p2_reverse_7937_comb[14:0] == 15'h0000, p2_reverse_7937_comb[14] && p2_reverse_7937_comb[13:0] == 14'h0000, p2_reverse_7937_comb[13] && p2_reverse_7937_comb[12:0] == 13'h0000, p2_reverse_7937_comb[12] && p2_reverse_7937_comb[11:0] == 12'h000, p2_reverse_7937_comb[11] && p2_reverse_7937_comb[10:0] == 11'h000, p2_reverse_7937_comb[10] && p2_reverse_7937_comb[9:0] == 10'h000, p2_reverse_7937_comb[9] && p2_reverse_7937_comb[8:0] == 9'h000, p2_reverse_7937_comb[8] && p2_reverse_7937_comb[7:0] == 8'h00, p2_reverse_7937_comb[7] && p2_reverse_7937_comb[6:0] == 7'h00, p2_reverse_7937_comb[6] && p2_reverse_7937_comb[5:0] == 6'h00, p2_reverse_7937_comb[5] && p2_reverse_7937_comb[4:0] == 5'h00, p2_reverse_7937_comb[4] && p2_reverse_7937_comb[3:0] == 4'h0, p2_reverse_7937_comb[3] && p2_reverse_7937_comb[2:0] == 3'h0, p2_reverse_7937_comb[2] && p2_reverse_7937_comb[1:0] == 2'h0, p2_reverse_7937_comb[1] && !p2_reverse_7937_comb[0], p2_reverse_7937_comb[0]};
  assign p2_one_hot_7940_comb = {p2_reverse_7938_comb[27:0] == 28'h000_0000, p2_reverse_7938_comb[27] && p2_reverse_7938_comb[26:0] == 27'h000_0000, p2_reverse_7938_comb[26] && p2_reverse_7938_comb[25:0] == 26'h000_0000, p2_reverse_7938_comb[25] && p2_reverse_7938_comb[24:0] == 25'h000_0000, p2_reverse_7938_comb[24] && p2_reverse_7938_comb[23:0] == 24'h00_0000, p2_reverse_7938_comb[23] && p2_reverse_7938_comb[22:0] == 23'h00_0000, p2_reverse_7938_comb[22] && p2_reverse_7938_comb[21:0] == 22'h00_0000, p2_reverse_7938_comb[21] && p2_reverse_7938_comb[20:0] == 21'h00_0000, p2_reverse_7938_comb[20] && p2_reverse_7938_comb[19:0] == 20'h0_0000, p2_reverse_7938_comb[19] && p2_reverse_7938_comb[18:0] == 19'h0_0000, p2_reverse_7938_comb[18] && p2_reverse_7938_comb[17:0] == 18'h0_0000, p2_reverse_7938_comb[17] && p2_reverse_7938_comb[16:0] == 17'h0_0000, p2_reverse_7938_comb[16] && p2_reverse_7938_comb[15:0] == 16'h0000, p2_reverse_7938_comb[15] && p2_reverse_7938_comb[14:0] == 15'h0000, p2_reverse_7938_comb[14] && p2_reverse_7938_comb[13:0] == 14'h0000, p2_reverse_7938_comb[13] && p2_reverse_7938_comb[12:0] == 13'h0000, p2_reverse_7938_comb[12] && p2_reverse_7938_comb[11:0] == 12'h000, p2_reverse_7938_comb[11] && p2_reverse_7938_comb[10:0] == 11'h000, p2_reverse_7938_comb[10] && p2_reverse_7938_comb[9:0] == 10'h000, p2_reverse_7938_comb[9] && p2_reverse_7938_comb[8:0] == 9'h000, p2_reverse_7938_comb[8] && p2_reverse_7938_comb[7:0] == 8'h00, p2_reverse_7938_comb[7] && p2_reverse_7938_comb[6:0] == 7'h00, p2_reverse_7938_comb[6] && p2_reverse_7938_comb[5:0] == 6'h00, p2_reverse_7938_comb[5] && p2_reverse_7938_comb[4:0] == 5'h00, p2_reverse_7938_comb[4] && p2_reverse_7938_comb[3:0] == 4'h0, p2_reverse_7938_comb[3] && p2_reverse_7938_comb[2:0] == 3'h0, p2_reverse_7938_comb[2] && p2_reverse_7938_comb[1:0] == 2'h0, p2_reverse_7938_comb[1] && !p2_reverse_7938_comb[0], p2_reverse_7938_comb[0]};
  assign p2_encode_7941_comb = {p2_one_hot_7939_comb[16] | p2_one_hot_7939_comb[17] | p2_one_hot_7939_comb[18] | p2_one_hot_7939_comb[19] | p2_one_hot_7939_comb[20] | p2_one_hot_7939_comb[21] | p2_one_hot_7939_comb[22] | p2_one_hot_7939_comb[23] | p2_one_hot_7939_comb[24] | p2_one_hot_7939_comb[25] | p2_one_hot_7939_comb[26] | p2_one_hot_7939_comb[27] | p2_one_hot_7939_comb[28], p2_one_hot_7939_comb[8] | p2_one_hot_7939_comb[9] | p2_one_hot_7939_comb[10] | p2_one_hot_7939_comb[11] | p2_one_hot_7939_comb[12] | p2_one_hot_7939_comb[13] | p2_one_hot_7939_comb[14] | p2_one_hot_7939_comb[15] | p2_one_hot_7939_comb[24] | p2_one_hot_7939_comb[25] | p2_one_hot_7939_comb[26] | p2_one_hot_7939_comb[27] | p2_one_hot_7939_comb[28], p2_one_hot_7939_comb[4] | p2_one_hot_7939_comb[5] | p2_one_hot_7939_comb[6] | p2_one_hot_7939_comb[7] | p2_one_hot_7939_comb[12] | p2_one_hot_7939_comb[13] | p2_one_hot_7939_comb[14] | p2_one_hot_7939_comb[15] | p2_one_hot_7939_comb[20] | p2_one_hot_7939_comb[21] | p2_one_hot_7939_comb[22] | p2_one_hot_7939_comb[23] | p2_one_hot_7939_comb[28], p2_one_hot_7939_comb[2] | p2_one_hot_7939_comb[3] | p2_one_hot_7939_comb[6] | p2_one_hot_7939_comb[7] | p2_one_hot_7939_comb[10] | p2_one_hot_7939_comb[11] | p2_one_hot_7939_comb[14] | p2_one_hot_7939_comb[15] | p2_one_hot_7939_comb[18] | p2_one_hot_7939_comb[19] | p2_one_hot_7939_comb[22] | p2_one_hot_7939_comb[23] | p2_one_hot_7939_comb[26] | p2_one_hot_7939_comb[27], p2_one_hot_7939_comb[1] | p2_one_hot_7939_comb[3] | p2_one_hot_7939_comb[5] | p2_one_hot_7939_comb[7] | p2_one_hot_7939_comb[9] | p2_one_hot_7939_comb[11] | p2_one_hot_7939_comb[13] | p2_one_hot_7939_comb[15] | p2_one_hot_7939_comb[17] | p2_one_hot_7939_comb[19] | p2_one_hot_7939_comb[21] | p2_one_hot_7939_comb[23] | p2_one_hot_7939_comb[25] | p2_one_hot_7939_comb[27]};
  assign p2_encode_7942_comb = {p2_one_hot_7940_comb[16] | p2_one_hot_7940_comb[17] | p2_one_hot_7940_comb[18] | p2_one_hot_7940_comb[19] | p2_one_hot_7940_comb[20] | p2_one_hot_7940_comb[21] | p2_one_hot_7940_comb[22] | p2_one_hot_7940_comb[23] | p2_one_hot_7940_comb[24] | p2_one_hot_7940_comb[25] | p2_one_hot_7940_comb[26] | p2_one_hot_7940_comb[27] | p2_one_hot_7940_comb[28], p2_one_hot_7940_comb[8] | p2_one_hot_7940_comb[9] | p2_one_hot_7940_comb[10] | p2_one_hot_7940_comb[11] | p2_one_hot_7940_comb[12] | p2_one_hot_7940_comb[13] | p2_one_hot_7940_comb[14] | p2_one_hot_7940_comb[15] | p2_one_hot_7940_comb[24] | p2_one_hot_7940_comb[25] | p2_one_hot_7940_comb[26] | p2_one_hot_7940_comb[27] | p2_one_hot_7940_comb[28], p2_one_hot_7940_comb[4] | p2_one_hot_7940_comb[5] | p2_one_hot_7940_comb[6] | p2_one_hot_7940_comb[7] | p2_one_hot_7940_comb[12] | p2_one_hot_7940_comb[13] | p2_one_hot_7940_comb[14] | p2_one_hot_7940_comb[15] | p2_one_hot_7940_comb[20] | p2_one_hot_7940_comb[21] | p2_one_hot_7940_comb[22] | p2_one_hot_7940_comb[23] | p2_one_hot_7940_comb[28], p2_one_hot_7940_comb[2] | p2_one_hot_7940_comb[3] | p2_one_hot_7940_comb[6] | p2_one_hot_7940_comb[7] | p2_one_hot_7940_comb[10] | p2_one_hot_7940_comb[11] | p2_one_hot_7940_comb[14] | p2_one_hot_7940_comb[15] | p2_one_hot_7940_comb[18] | p2_one_hot_7940_comb[19] | p2_one_hot_7940_comb[22] | p2_one_hot_7940_comb[23] | p2_one_hot_7940_comb[26] | p2_one_hot_7940_comb[27], p2_one_hot_7940_comb[1] | p2_one_hot_7940_comb[3] | p2_one_hot_7940_comb[5] | p2_one_hot_7940_comb[7] | p2_one_hot_7940_comb[9] | p2_one_hot_7940_comb[11] | p2_one_hot_7940_comb[13] | p2_one_hot_7940_comb[15] | p2_one_hot_7940_comb[17] | p2_one_hot_7940_comb[19] | p2_one_hot_7940_comb[21] | p2_one_hot_7940_comb[23] | p2_one_hot_7940_comb[25] | p2_one_hot_7940_comb[27]};
  assign p2_carry_bit_comb = p2_abs_fraction_comb[27];
  assign p2_cancel_comb = p2_encode_7941_comb[1] | p2_encode_7941_comb[2] | p2_encode_7941_comb[3] | p2_encode_7941_comb[4];
  assign p2_carry_bit__1_comb = p2_abs_fraction__1_comb[27];
  assign p2_cancel__1_comb = p2_encode_7942_comb[1] | p2_encode_7942_comb[2] | p2_encode_7942_comb[3] | p2_encode_7942_comb[4];
  assign p2_leading_zeroes_comb = {23'h00_0000, p2_encode_7941_comb};
  assign p2_leading_zeroes__1_comb = {23'h00_0000, p2_encode_7942_comb};
  assign p2_and_7969_comb = ~p2_carry_bit_comb & ~p2_cancel_comb;
  assign p2_and_7970_comb = ~p2_carry_bit_comb & p2_cancel_comb;
  assign p2_and_7971_comb = p2_carry_bit_comb & ~p2_cancel_comb;
  assign p2_carry_fraction_comb = p2_abs_fraction_comb[27:1];
  assign p2_add_7975_comb = p2_leading_zeroes_comb + 28'hfff_ffff;
  assign p2_and_7976_comb = ~p2_carry_bit__1_comb & ~p2_cancel__1_comb;
  assign p2_and_7977_comb = ~p2_carry_bit__1_comb & p2_cancel__1_comb;
  assign p2_and_7978_comb = p2_carry_bit__1_comb & ~p2_cancel__1_comb;
  assign p2_carry_fraction__2_comb = p2_abs_fraction__1_comb[27:1];
  assign p2_add_7982_comb = p2_leading_zeroes__1_comb + 28'hfff_ffff;
  assign p2_concat_7983_comb = {p2_and_7969_comb, p2_and_7970_comb, p2_and_7971_comb};
  assign p2_carry_fraction__1_comb = p2_carry_fraction_comb | {26'h000_0000, p2_abs_fraction_comb[0]};
  assign p2_cancel_fraction_comb = p2_add_7975_comb >= 28'h000_001b ? 27'h000_0000 : p2_abs_fraction_comb[26:0] << p2_add_7975_comb;
  assign p2_concat_7986_comb = {p2_and_7976_comb, p2_and_7977_comb, p2_and_7978_comb};
  assign p2_carry_fraction__3_comb = p2_carry_fraction__2_comb | {26'h000_0000, p2_abs_fraction__1_comb[0]};
  assign p2_cancel_fraction__1_comb = p2_add_7982_comb >= 28'h000_001b ? 27'h000_0000 : p2_abs_fraction__1_comb[26:0] << p2_add_7982_comb;
  assign p2_shifted_fraction_comb = p2_carry_fraction__1_comb & {27{p2_concat_7983_comb[0]}} | p2_cancel_fraction_comb & {27{p2_concat_7983_comb[1]}} | p2_abs_fraction_comb[26:0] & {27{p2_concat_7983_comb[2]}};
  assign p2_shifted_fraction__1_comb = p2_carry_fraction__3_comb & {27{p2_concat_7986_comb[0]}} | p2_cancel_fraction__1_comb & {27{p2_concat_7986_comb[1]}} | p2_abs_fraction__1_comb[26:0] & {27{p2_concat_7986_comb[2]}};
  assign p2_normal_chunk_comb = p2_shifted_fraction_comb[2:0];
  assign p2_half_way_chunk_comb = p2_shifted_fraction_comb[3:2];
  assign p2_normal_chunk__1_comb = p2_shifted_fraction__1_comb[2:0];
  assign p2_half_way_chunk__1_comb = p2_shifted_fraction__1_comb[3:2];
  assign p2_add_8010_comb = {1'h0, p2_shifted_fraction_comb[26:3]} + 25'h000_0001;
  assign p2_add_8014_comb = {1'h0, p2_shifted_fraction__1_comb[26:3]} + 25'h000_0001;
  assign p2_do_round_up__5_comb = p2_normal_chunk_comb > 3'h4 | p2_half_way_chunk_comb == 2'h3;
  assign p2_do_round_up__6_comb = p2_normal_chunk__1_comb > 3'h4 | p2_half_way_chunk__1_comb == 2'h3;
  assign p2_rounded_fraction_comb = p2_do_round_up__5_comb ? {p2_add_8010_comb, p2_normal_chunk_comb} : {1'h0, p2_shifted_fraction_comb};
  assign p2_rounded_fraction__1_comb = p2_do_round_up__6_comb ? {p2_add_8014_comb, p2_normal_chunk__1_comb} : {1'h0, p2_shifted_fraction__1_comb};
  assign p2_rounding_carry_comb = p2_rounded_fraction_comb[27];
  assign p2_rounding_carry__1_comb = p2_rounded_fraction__1_comb[27];
  assign p2_add_8034_comb = {1'h0, p1_greater_exp_bexp} + {8'h00, p2_rounding_carry_comb};
  assign p2_add_8036_comb = {1'h0, p1_greater_exp_bexp__1} + {8'h00, p2_rounding_carry__1_comb};
  assign p2_add_8043_comb = {1'h0, p2_add_8034_comb} + 10'h001;
  assign p2_add_8045_comb = {1'h0, p2_add_8036_comb} + 10'h001;
  assign p2_wide_exponent_comb = p2_add_8043_comb - {5'h00, p2_encode_7941_comb};
  assign p2_wide_exponent__3_comb = p2_add_8045_comb - {5'h00, p2_encode_7942_comb};
  assign p2_wide_exponent__1_comb = p2_wide_exponent_comb & {10{p1_ne_7808}};
  assign p2_wide_exponent__4_comb = p2_wide_exponent__3_comb & {10{p1_ne_7809}};
  assign p2_wide_exponent__2_comb = p2_wide_exponent__1_comb[8:0] & {9{~p2_wide_exponent__1_comb[9]}};
  assign p2_wide_exponent__5_comb = p2_wide_exponent__4_comb[8:0] & {9{~p2_wide_exponent__4_comb[9]}};
  assign p2_add_8089_comb = {2'h0, p2_rounding_carry_comb} + 3'h3;
  assign p2_add_8092_comb = {2'h0, p2_rounding_carry__1_comb} + 3'h3;
  assign p2_shrl_8095_comb = p2_rounded_fraction_comb >> p2_add_8089_comb;
  assign p2_nor_8097_comb = ~(p2_wide_exponent__2_comb[8] | p2_wide_exponent__2_comb[0] & p2_wide_exponent__2_comb[1] & p2_wide_exponent__2_comb[2] & p2_wide_exponent__2_comb[3] & p2_wide_exponent__2_comb[4] & p2_wide_exponent__2_comb[5] & p2_wide_exponent__2_comb[6] & p2_wide_exponent__2_comb[7]);
  assign p2_shrl_8098_comb = p2_rounded_fraction__1_comb >> p2_add_8092_comb;
  assign p2_nor_8100_comb = ~(p2_wide_exponent__5_comb[8] | p2_wide_exponent__5_comb[0] & p2_wide_exponent__5_comb[1] & p2_wide_exponent__5_comb[2] & p2_wide_exponent__5_comb[3] & p2_wide_exponent__5_comb[4] & p2_wide_exponent__5_comb[5] & p2_wide_exponent__5_comb[6] & p2_wide_exponent__5_comb[7]);
  assign p2_result_fraction__13_comb = p2_shrl_8095_comb[22:0];
  assign p2_result_fraction__15_comb = p2_shrl_8098_comb[22:0];
  assign p2_result_fraction__14_comb = p2_result_fraction__13_comb & {23{~(~(p2_wide_exponent__2_comb[1] | p2_wide_exponent__2_comb[2] | p2_wide_exponent__2_comb[3] | p2_wide_exponent__2_comb[4] | p2_wide_exponent__2_comb[5] | p2_wide_exponent__2_comb[6] | p2_wide_exponent__2_comb[7] | p2_wide_exponent__2_comb[8] | p2_wide_exponent__2_comb[0]))}} & {23{p2_nor_8097_comb}} & {23{p1_nor_7854}};
  assign p2_nan_fraction__14_comb = 23'h40_0000;
  assign p2_high_exp__36_comb = 8'hff;
  assign p2_result_fraction__16_comb = p2_result_fraction__15_comb & {23{~(~(p2_wide_exponent__5_comb[1] | p2_wide_exponent__5_comb[2] | p2_wide_exponent__5_comb[3] | p2_wide_exponent__5_comb[4] | p2_wide_exponent__5_comb[5] | p2_wide_exponent__5_comb[6] | p2_wide_exponent__5_comb[7] | p2_wide_exponent__5_comb[8] | p2_wide_exponent__5_comb[0]))}} & {23{p2_nor_8100_comb}} & {23{p1_nor_7858}};
  assign p2_nan_fraction__15_comb = 23'h40_0000;
  assign p2_high_exp__37_comb = 8'hff;
  assign p2_result_fraction__17_comb = p1_is_result_nan__5 ? p2_nan_fraction__14_comb : p2_result_fraction__14_comb;
  assign p2_result_exponent__2_comb = p1_is_result_nan__5 | p1_is_operand_inf | ~p2_nor_8097_comb ? p2_high_exp__36_comb : p2_wide_exponent__2_comb[7:0];
  assign p2_result_fraction__18_comb = p1_is_result_nan__6 ? p2_nan_fraction__15_comb : p2_result_fraction__16_comb;
  assign p2_result_exponent__1_comb = p1_is_result_nan__6 | p1_is_operand_inf__1 | ~p2_nor_8100_comb ? p2_high_exp__37_comb : p2_wide_exponent__5_comb[7:0];
  assign p2_add_8152_comb = p1_in0_r_bexp__6[7:2] + 6'h07;
  assign p2_ugt_8154_comb = p1_in0_r_bexp__6 > p2_result_exponent__2_comb;
  assign p2_add_8163_comb = p1_in0_i_bexp__6[7:2] + 6'h07;
  assign p2_ugt_8165_comb = p1_in0_i_bexp__6 > p2_result_exponent__1_comb;
  assign p2_result_sign__9_comb = ~(~p1_bit_slice_7804 | p1_greater_exp_sign) | ~(p1_bit_slice_7804 | p1_fraction_is_zero | ~p1_greater_exp_sign);
  assign p2_result_sign__11_comb = ~(~p1_bit_slice_7805 | p1_greater_exp_sign__1) | ~(p1_bit_slice_7805 | p1_fraction_is_zero__1 | ~p1_greater_exp_sign__1);
  assign p2_add_8158_comb = p2_result_exponent__2_comb[7:2] + 6'h07;
  assign p2_add_8169_comb = p2_result_exponent__1_comb[7:2] + 6'h07;
  assign p2_wide_x__4_comb = {{2'h0, p1_in0_r_fraction__6} | 25'h080_0000, 3'h0};
  assign p2_greater_exp_bexp__2_comb = p2_ugt_8154_comb ? p1_in0_r_bexp__6 : p2_result_exponent__2_comb;
  assign p2_wide_x__6_comb = {{2'h0, p1_in0_i_fraction__6} | 25'h080_0000, 3'h0};
  assign p2_greater_exp_bexp__3_comb = p2_ugt_8165_comb ? p1_in0_i_bexp__6 : p2_result_exponent__1_comb;
  assign p2_high_exp__39_comb = 8'hff;
  assign p2_result_sign__10_comb = p1_is_operand_inf ? p1_not_7874 : p2_result_sign__9_comb;
  assign p2_high_exp__41_comb = 8'hff;
  assign p2_result_sign__12_comb = p1_is_operand_inf__1 ? p1_not_7875 : p2_result_sign__11_comb;
  assign p2_wide_y__4_comb = {{2'h0, p2_result_fraction__17_comb} | 25'h080_0000, 3'h0};
  assign p2_wide_y__6_comb = {{2'h0, p2_result_fraction__18_comb} | 25'h080_0000, 3'h0};
  assign p2_wide_x__5_comb = p2_wide_x__4_comb & {28{p1_in0_r_bexp__6 != 8'h00}};
  assign p2_sub_8190_comb = {p2_add_8152_comb, p1_in0_r_bexp__6[1:0]} - p2_greater_exp_bexp__2_comb;
  assign p2_wide_x__7_comb = p2_wide_x__6_comb & {28{p1_in0_i_bexp__6 != 8'h00}};
  assign p2_sub_8194_comb = {p2_add_8163_comb, p1_in0_i_bexp__6[1:0]} - p2_greater_exp_bexp__3_comb;
  assign p2_high_exp__46_comb = 8'hff;
  assign p2_eq_8251_comb = p2_result_exponent__2_comb == p2_high_exp__39_comb;
  assign p2_eq_8252_comb = p2_result_fraction__17_comb == 23'h00_0000;
  assign p2_high_exp__38_comb = 8'hff;
  assign p2_result_sign__13_comb = ~p1_is_result_nan__5 & p2_result_sign__10_comb;
  assign p2_high_exp__47_comb = 8'hff;
  assign p2_eq_8257_comb = p2_result_exponent__1_comb == p2_high_exp__41_comb;
  assign p2_eq_8258_comb = p2_result_fraction__18_comb == 23'h00_0000;
  assign p2_high_exp__40_comb = 8'hff;
  assign p2_result_sign__14_comb = ~p1_is_result_nan__6 & p2_result_sign__12_comb;
  assign p2_wide_y__5_comb = p2_wide_y__4_comb & {28{p2_result_exponent__2_comb != 8'h00}};
  assign p2_sub_8192_comb = {p2_add_8158_comb, p2_result_exponent__2_comb[1:0]} - p2_greater_exp_bexp__2_comb;
  assign p2_wide_y__7_comb = p2_wide_y__6_comb & {28{p2_result_exponent__1_comb != 8'h00}};
  assign p2_sub_8196_comb = {p2_add_8169_comb, p2_result_exponent__1_comb[1:0]} - p2_greater_exp_bexp__3_comb;
  assign p2_dropped_x__2_comb = p2_sub_8190_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__5_comb << p2_sub_8190_comb;
  assign p2_dropped_x__3_comb = p2_sub_8194_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__7_comb << p2_sub_8194_comb;
  assign p2_ne_8262_comb = p1_in0_r_fraction__6 != 23'h00_0000;
  assign p2_nand_8263_comb = ~(p2_eq_8251_comb & p2_eq_8252_comb);
  assign p2_eq_8264_comb = p1_in0_r_bexp__6 == p2_high_exp__38_comb;
  assign p2_eq_8265_comb = p1_in0_r_fraction__6 == 23'h00_0000;
  assign p2_re__1_sign_comb = ~p2_result_sign__13_comb;
  assign p2_ne_8267_comb = p1_in0_i_fraction__6 != 23'h00_0000;
  assign p2_nand_8268_comb = ~(p2_eq_8257_comb & p2_eq_8258_comb);
  assign p2_eq_8269_comb = p1_in0_i_bexp__6 == p2_high_exp__40_comb;
  assign p2_eq_8270_comb = p1_in0_i_fraction__6 == 23'h00_0000;
  assign p2_im__1_sign_comb = ~p2_result_sign__14_comb;
  assign p2_dropped_y__2_comb = p2_sub_8192_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__5_comb << p2_sub_8192_comb;
  assign p2_dropped_y__3_comb = p2_sub_8196_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__7_comb << p2_sub_8196_comb;
  assign p2_nor_8272_comb = ~(p1_in0_r_bexp__6 != p2_high_exp__46_comb | p2_ne_8262_comb | p1_in0_r_sign__2);
  assign p2_nor_8273_comb = ~(p2_nand_8263_comb | p2_result_sign__13_comb);
  assign p2_and_8274_comb = p2_eq_8264_comb & p2_eq_8265_comb & p1_in0_r_sign__2;
  assign p2_nor_8275_comb = ~(p2_nand_8263_comb | p2_re__1_sign_comb);
  assign p2_nor_8277_comb = ~(p1_in0_i_bexp__6 != p2_high_exp__47_comb | p2_ne_8267_comb | p1_in0_i_sign__2);
  assign p2_nor_8278_comb = ~(p2_nand_8268_comb | p2_result_sign__14_comb);
  assign p2_and_8279_comb = p2_eq_8269_comb & p2_eq_8270_comb & p1_in0_i_sign__2;
  assign p2_nor_8280_comb = ~(p2_nand_8268_comb | p2_im__1_sign_comb);
  assign p2_shift_x__2_comb = p2_greater_exp_bexp__2_comb - p1_in0_r_bexp__6;
  assign p2_sticky_x__2_comb = p2_dropped_x__2_comb[27:3] != 25'h000_0000;
  assign p2_shift_x__3_comb = p2_greater_exp_bexp__3_comb - p1_in0_i_bexp__6;
  assign p2_sticky_x__3_comb = p2_dropped_x__3_comb[27:3] != 25'h000_0000;
  assign p2_has_pos_inf__2_comb = p2_nor_8272_comb | p2_nor_8273_comb;
  assign p2_has_neg_inf__2_comb = p2_and_8274_comb | p2_nor_8275_comb;
  assign p2_has_pos_inf__3_comb = p2_nor_8277_comb | p2_nor_8278_comb;
  assign p2_has_neg_inf__3_comb = p2_and_8279_comb | p2_nor_8280_comb;
  assign p2_has_pos_inf__4_comb = p2_nor_8272_comb | p2_nor_8275_comb;
  assign p2_has_neg_inf__4_comb = p2_and_8274_comb | p2_nor_8273_comb;
  assign p2_has_pos_inf__5_comb = p2_nor_8277_comb | p2_nor_8280_comb;
  assign p2_has_neg_inf__5_comb = p2_and_8279_comb | p2_nor_8278_comb;
  assign p2_shift_y__2_comb = p2_greater_exp_bexp__2_comb - p2_result_exponent__2_comb;
  assign p2_sticky_y__2_comb = p2_dropped_y__2_comb[27:3] != 25'h000_0000;
  assign p2_shift_y__3_comb = p2_greater_exp_bexp__3_comb - p2_result_exponent__1_comb;
  assign p2_sticky_y__3_comb = p2_dropped_y__3_comb[27:3] != 25'h000_0000;
  assign p2_shifted_x__2_comb = p2_shift_x__2_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__5_comb >> p2_shift_x__2_comb;
  assign p2_shifted_x__3_comb = p2_shift_x__3_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__7_comb >> p2_shift_x__3_comb;
  assign p2_and_8284_comb = p2_eq_8264_comb & p2_eq_8265_comb;
  assign p2_and_8285_comb = p2_eq_8251_comb & p2_eq_8252_comb;
  assign p2_and_8289_comb = p2_eq_8269_comb & p2_eq_8270_comb;
  assign p2_and_8290_comb = p2_eq_8257_comb & p2_eq_8258_comb;
  assign p2_and_8295_comb = p2_eq_8264_comb & p2_ne_8262_comb;
  assign p2_and_8296_comb = p2_eq_8251_comb & p2_result_fraction__17_comb != 23'h00_0000;
  assign p2_and_8299_comb = p2_eq_8269_comb & p2_ne_8267_comb;
  assign p2_and_8300_comb = p2_eq_8257_comb & p2_result_fraction__18_comb != 23'h00_0000;
  assign p2_shifted_y__2_comb = p2_shift_y__2_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__5_comb >> p2_shift_y__2_comb;
  assign p2_concat_8236_comb = {27'h000_0000, p2_sticky_y__2_comb};
  assign p2_shifted_y__3_comb = p2_shift_y__3_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__7_comb >> p2_shift_y__3_comb;
  assign p2_concat_8240_comb = {27'h000_0000, p2_sticky_y__3_comb};
  assign p2_addend_x__4_comb = p2_shifted_x__2_comb | {27'h000_0000, p2_sticky_x__2_comb};
  assign p2_addend_x__6_comb = p2_shifted_x__3_comb | {27'h000_0000, p2_sticky_x__3_comb};
  assign p2_nor_8298_comb = ~(p2_and_8284_comb | p2_and_8285_comb);
  assign p2_nor_8302_comb = ~(p2_and_8289_comb | p2_and_8290_comb);
  assign p2_is_result_nan__7_comb = p2_and_8295_comb | p2_and_8296_comb | p2_has_pos_inf__2_comb & p2_has_neg_inf__2_comb;
  assign p2_is_operand_inf__2_comb = p2_and_8284_comb | p2_and_8285_comb;
  assign p2_not_8307_comb = ~p2_has_pos_inf__2_comb;
  assign p2_is_result_nan__8_comb = p2_and_8299_comb | p2_and_8300_comb | p2_has_pos_inf__3_comb & p2_has_neg_inf__3_comb;
  assign p2_is_operand_inf__3_comb = p2_and_8289_comb | p2_and_8290_comb;
  assign p2_not_8310_comb = ~p2_has_pos_inf__3_comb;
  assign p2_is_result_nan__9_comb = p2_and_8295_comb | p2_and_8296_comb | p2_has_pos_inf__4_comb & p2_has_neg_inf__4_comb;
  assign p2_not_8312_comb = ~p2_has_pos_inf__4_comb;
  assign p2_is_result_nan__10_comb = p2_and_8299_comb | p2_and_8300_comb | p2_has_pos_inf__5_comb & p2_has_neg_inf__5_comb;
  assign p2_not_8314_comb = ~p2_has_pos_inf__5_comb;

  // Registers for pipe stage 2:
  reg p2_ugt_8154;
  reg p2_ugt_8165;
  reg [7:0] p2_greater_exp_bexp__2;
  reg [7:0] p2_greater_exp_bexp__3;
  reg p2_result_sign__13;
  reg p2_result_sign__14;
  reg p2_in0_r_sign__2;
  reg [27:0] p2_shifted_y__2;
  reg [27:0] p2_concat_8236;
  reg p2_in0_i_sign__2;
  reg [27:0] p2_shifted_y__3;
  reg [27:0] p2_concat_8240;
  reg p2_re__1_sign;
  reg p2_im__1_sign;
  reg [27:0] p2_addend_x__4;
  reg [27:0] p2_addend_x__6;
  reg p2_nor_8298;
  reg p2_nor_8302;
  reg p2_is_result_nan__7;
  reg p2_is_operand_inf__2;
  reg p2_not_8307;
  reg p2_is_result_nan__8;
  reg p2_is_operand_inf__3;
  reg p2_not_8310;
  reg p2_is_result_nan__9;
  reg p2_not_8312;
  reg p2_is_result_nan__10;
  reg p2_not_8314;
  always_ff @ (posedge clk) begin
    p2_ugt_8154 <= p2_ugt_8154_comb;
    p2_ugt_8165 <= p2_ugt_8165_comb;
    p2_greater_exp_bexp__2 <= p2_greater_exp_bexp__2_comb;
    p2_greater_exp_bexp__3 <= p2_greater_exp_bexp__3_comb;
    p2_result_sign__13 <= p2_result_sign__13_comb;
    p2_result_sign__14 <= p2_result_sign__14_comb;
    p2_in0_r_sign__2 <= p1_in0_r_sign__2;
    p2_shifted_y__2 <= p2_shifted_y__2_comb;
    p2_concat_8236 <= p2_concat_8236_comb;
    p2_in0_i_sign__2 <= p1_in0_i_sign__2;
    p2_shifted_y__3 <= p2_shifted_y__3_comb;
    p2_concat_8240 <= p2_concat_8240_comb;
    p2_re__1_sign <= p2_re__1_sign_comb;
    p2_im__1_sign <= p2_im__1_sign_comb;
    p2_addend_x__4 <= p2_addend_x__4_comb;
    p2_addend_x__6 <= p2_addend_x__6_comb;
    p2_nor_8298 <= p2_nor_8298_comb;
    p2_nor_8302 <= p2_nor_8302_comb;
    p2_is_result_nan__7 <= p2_is_result_nan__7_comb;
    p2_is_operand_inf__2 <= p2_is_operand_inf__2_comb;
    p2_not_8307 <= p2_not_8307_comb;
    p2_is_result_nan__8 <= p2_is_result_nan__8_comb;
    p2_is_operand_inf__3 <= p2_is_operand_inf__3_comb;
    p2_not_8310 <= p2_not_8310_comb;
    p2_is_result_nan__9 <= p2_is_result_nan__9_comb;
    p2_not_8312 <= p2_not_8312_comb;
    p2_is_result_nan__10 <= p2_is_result_nan__10_comb;
    p2_not_8314 <= p2_not_8314_comb;
  end

  // ===== Pipe stage 3:
  wire p3_greater_exp_sign__2_comb;
  wire [27:0] p3_addend_y__4_comb;
  wire p3_greater_exp_sign__3_comb;
  wire [27:0] p3_addend_y__6_comb;
  wire p3_greater_exp_sign__4_comb;
  wire p3_greater_exp_sign__5_comb;
  wire [27:0] p3_addend_x__5_comb;
  wire [27:0] p3_addend_y__5_comb;
  wire [27:0] p3_addend_x__7_comb;
  wire [27:0] p3_addend_y__7_comb;
  wire [27:0] p3_addend_x__9_comb;
  wire [27:0] p3_addend_y__9_comb;
  wire [27:0] p3_addend_x__11_comb;
  wire [27:0] p3_addend_y__11_comb;
  wire [28:0] p3_fraction__35_comb;
  wire [28:0] p3_fraction__36_comb;
  wire [28:0] p3_fraction__37_comb;
  wire [28:0] p3_fraction__38_comb;
  wire [27:0] p3_abs_fraction__2_comb;
  wire [27:0] p3_abs_fraction__3_comb;
  wire [27:0] p3_abs_fraction__4_comb;
  wire [27:0] p3_abs_fraction__5_comb;
  wire [27:0] p3_reverse_8431_comb;
  wire [27:0] p3_reverse_8432_comb;
  wire [27:0] p3_reverse_8433_comb;
  wire [27:0] p3_reverse_8434_comb;
  wire [28:0] p3_one_hot_8435_comb;
  wire [28:0] p3_one_hot_8436_comb;
  wire [28:0] p3_one_hot_8437_comb;
  wire [28:0] p3_one_hot_8438_comb;
  wire [4:0] p3_encode_8439_comb;
  wire [4:0] p3_encode_8440_comb;
  wire [4:0] p3_encode_8441_comb;
  wire [4:0] p3_encode_8442_comb;
  wire p3_carry_bit__2_comb;
  wire p3_cancel__2_comb;
  wire p3_carry_bit__3_comb;
  wire p3_cancel__3_comb;
  wire p3_carry_bit__4_comb;
  wire p3_cancel__4_comb;
  wire p3_carry_bit__5_comb;
  wire p3_cancel__5_comb;
  wire [27:0] p3_leading_zeroes__2_comb;
  wire [27:0] p3_leading_zeroes__3_comb;
  wire [27:0] p3_leading_zeroes__4_comb;
  wire [27:0] p3_leading_zeroes__5_comb;
  wire p3_and_8495_comb;
  wire p3_and_8496_comb;
  wire p3_and_8497_comb;
  wire [26:0] p3_carry_fraction__4_comb;
  wire [27:0] p3_add_8501_comb;
  wire p3_and_8502_comb;
  wire p3_and_8503_comb;
  wire p3_and_8504_comb;
  wire [26:0] p3_carry_fraction__6_comb;
  wire [27:0] p3_add_8508_comb;
  wire p3_and_8509_comb;
  wire p3_and_8510_comb;
  wire p3_and_8511_comb;
  wire [26:0] p3_carry_fraction__8_comb;
  wire [27:0] p3_add_8515_comb;
  wire p3_and_8516_comb;
  wire p3_and_8517_comb;
  wire p3_and_8518_comb;
  wire [26:0] p3_carry_fraction__10_comb;
  wire [27:0] p3_add_8522_comb;
  wire [2:0] p3_concat_8523_comb;
  wire [26:0] p3_carry_fraction__5_comb;
  wire [26:0] p3_cancel_fraction__2_comb;
  wire [2:0] p3_concat_8526_comb;
  wire [26:0] p3_carry_fraction__7_comb;
  wire [26:0] p3_cancel_fraction__3_comb;
  wire [2:0] p3_concat_8529_comb;
  wire [26:0] p3_carry_fraction__9_comb;
  wire [26:0] p3_cancel_fraction__4_comb;
  wire [2:0] p3_concat_8532_comb;
  wire [26:0] p3_carry_fraction__11_comb;
  wire [26:0] p3_cancel_fraction__5_comb;
  wire [26:0] p3_shifted_fraction__2_comb;
  wire [26:0] p3_shifted_fraction__3_comb;
  wire [26:0] p3_shifted_fraction__4_comb;
  wire [26:0] p3_shifted_fraction__5_comb;
  wire [2:0] p3_normal_chunk__2_comb;
  wire [1:0] p3_half_way_chunk__2_comb;
  wire [2:0] p3_normal_chunk__3_comb;
  wire [1:0] p3_half_way_chunk__3_comb;
  wire [2:0] p3_normal_chunk__4_comb;
  wire [1:0] p3_half_way_chunk__4_comb;
  wire [2:0] p3_normal_chunk__5_comb;
  wire [1:0] p3_half_way_chunk__5_comb;
  wire [24:0] p3_add_8574_comb;
  wire [24:0] p3_add_8578_comb;
  wire [24:0] p3_add_8582_comb;
  wire [24:0] p3_add_8586_comb;
  wire p3_do_round_up__7_comb;
  wire p3_do_round_up__8_comb;
  wire p3_do_round_up__9_comb;
  wire p3_do_round_up__10_comb;
  wire [27:0] p3_rounded_fraction__2_comb;
  wire [27:0] p3_rounded_fraction__3_comb;
  wire [27:0] p3_rounded_fraction__4_comb;
  wire [27:0] p3_rounded_fraction__5_comb;
  wire p3_rounding_carry__2_comb;
  wire p3_rounding_carry__3_comb;
  wire p3_rounding_carry__4_comb;
  wire p3_rounding_carry__5_comb;
  wire [8:0] p3_concat_8613_comb;
  wire [8:0] p3_concat_8615_comb;
  wire [8:0] p3_add_8620_comb;
  wire [8:0] p3_add_8622_comb;
  wire [8:0] p3_add_8624_comb;
  wire [8:0] p3_add_8626_comb;
  wire [9:0] p3_add_8643_comb;
  wire [9:0] p3_add_8646_comb;
  wire [9:0] p3_add_8649_comb;
  wire [9:0] p3_add_8652_comb;
  wire [9:0] p3_wide_exponent__6_comb;
  wire [9:0] p3_wide_exponent__9_comb;
  wire [9:0] p3_wide_exponent__12_comb;
  wire [9:0] p3_wide_exponent__15_comb;
  wire [9:0] p3_wide_exponent__7_comb;
  wire [9:0] p3_wide_exponent__10_comb;
  wire [9:0] p3_wide_exponent__13_comb;
  wire [9:0] p3_wide_exponent__16_comb;
  wire [8:0] p3_wide_exponent__8_comb;
  wire [8:0] p3_wide_exponent__11_comb;
  wire [8:0] p3_wide_exponent__14_comb;
  wire [8:0] p3_wide_exponent__17_comb;
  wire p3_fraction_is_zero__2_comb;
  wire [2:0] p3_add_8747_comb;
  wire p3_fraction_is_zero__3_comb;
  wire [2:0] p3_add_8753_comb;
  wire p3_fraction_is_zero__4_comb;
  wire [2:0] p3_add_8759_comb;
  wire p3_fraction_is_zero__5_comb;
  wire [2:0] p3_add_8765_comb;
  wire p3_nor_8769_comb;
  wire [27:0] p3_shrl_8770_comb;
  wire p3_nor_8774_comb;
  wire [27:0] p3_shrl_8775_comb;
  wire p3_nor_8779_comb;
  wire [27:0] p3_shrl_8780_comb;
  wire p3_nor_8784_comb;
  wire [27:0] p3_shrl_8785_comb;
  wire p3_result_sign__15_comb;
  wire [22:0] p3_result_fraction__19_comb;
  wire [22:0] p3_sign_ext_8792_comb;
  wire p3_result_sign__17_comb;
  wire [22:0] p3_result_fraction__21_comb;
  wire [22:0] p3_sign_ext_8798_comb;
  wire p3_result_sign__20_comb;
  wire [22:0] p3_result_fraction__24_comb;
  wire p3_result_sign__23_comb;
  wire [22:0] p3_result_fraction__27_comb;
  wire p3_result_sign__16_comb;
  wire [7:0] p3_high_exp__42_comb;
  wire [22:0] p3_result_fraction__20_comb;
  wire [22:0] p3_nan_fraction__16_comb;
  wire p3_result_sign__18_comb;
  wire [7:0] p3_high_exp__43_comb;
  wire [22:0] p3_result_fraction__22_comb;
  wire [22:0] p3_nan_fraction__17_comb;
  wire p3_result_sign__21_comb;
  wire [7:0] p3_high_exp__44_comb;
  wire [22:0] p3_result_fraction__25_comb;
  wire [22:0] p3_nan_fraction__18_comb;
  wire p3_result_sign__24_comb;
  wire [7:0] p3_high_exp__45_comb;
  wire [22:0] p3_result_fraction__28_comb;
  wire [22:0] p3_nan_fraction__19_comb;
  wire p3_result_sign__19_comb;
  wire [7:0] p3_result_exponent__3_comb;
  wire [22:0] p3_result_fraction__23_comb;
  wire p3_result_sign__22_comb;
  wire [7:0] p3_result_exponent__4_comb;
  wire [22:0] p3_result_fraction__26_comb;
  wire p3_result_sign__25_comb;
  wire [7:0] p3_result_exponent__5_comb;
  wire [22:0] p3_result_fraction__29_comb;
  wire p3_result_sign__26_comb;
  wire [7:0] p3_result_exponent__6_comb;
  wire [22:0] p3_result_fraction__30_comb;
  wire [31:0] p3_out0_r_comb;
  wire [31:0] p3_out0_i_comb;
  wire [31:0] p3_out1_r_comb;
  wire [31:0] p3_out1_i_comb;
  wire [127:0] p3_tuple_8861_comb;
  assign p3_greater_exp_sign__2_comb = p2_ugt_8154 ? p2_in0_r_sign__2 : p2_result_sign__13;
  assign p3_addend_y__4_comb = p2_shifted_y__2 | p2_concat_8236;
  assign p3_greater_exp_sign__3_comb = p2_ugt_8165 ? p2_in0_i_sign__2 : p2_result_sign__14;
  assign p3_addend_y__6_comb = p2_shifted_y__3 | p2_concat_8240;
  assign p3_greater_exp_sign__4_comb = p2_ugt_8154 ? p2_in0_r_sign__2 : p2_re__1_sign;
  assign p3_greater_exp_sign__5_comb = p2_ugt_8165 ? p2_in0_i_sign__2 : p2_im__1_sign;
  assign p3_addend_x__5_comb = p2_in0_r_sign__2 ^ p3_greater_exp_sign__2_comb ? -p2_addend_x__4 : p2_addend_x__4;
  assign p3_addend_y__5_comb = p2_result_sign__13 ^ p3_greater_exp_sign__2_comb ? -p3_addend_y__4_comb : p3_addend_y__4_comb;
  assign p3_addend_x__7_comb = p2_in0_i_sign__2 ^ p3_greater_exp_sign__3_comb ? -p2_addend_x__6 : p2_addend_x__6;
  assign p3_addend_y__7_comb = p2_result_sign__14 ^ p3_greater_exp_sign__3_comb ? -p3_addend_y__6_comb : p3_addend_y__6_comb;
  assign p3_addend_x__9_comb = p2_in0_r_sign__2 ^ p3_greater_exp_sign__4_comb ? -p2_addend_x__4 : p2_addend_x__4;
  assign p3_addend_y__9_comb = p2_re__1_sign ^ p3_greater_exp_sign__4_comb ? -p3_addend_y__4_comb : p3_addend_y__4_comb;
  assign p3_addend_x__11_comb = p2_in0_i_sign__2 ^ p3_greater_exp_sign__5_comb ? -p2_addend_x__6 : p2_addend_x__6;
  assign p3_addend_y__11_comb = p2_im__1_sign ^ p3_greater_exp_sign__5_comb ? -p3_addend_y__6_comb : p3_addend_y__6_comb;
  assign p3_fraction__35_comb = {{1{p3_addend_x__5_comb[27]}}, p3_addend_x__5_comb} + {{1{p3_addend_y__5_comb[27]}}, p3_addend_y__5_comb};
  assign p3_fraction__36_comb = {{1{p3_addend_x__7_comb[27]}}, p3_addend_x__7_comb} + {{1{p3_addend_y__7_comb[27]}}, p3_addend_y__7_comb};
  assign p3_fraction__37_comb = {{1{p3_addend_x__9_comb[27]}}, p3_addend_x__9_comb} + {{1{p3_addend_y__9_comb[27]}}, p3_addend_y__9_comb};
  assign p3_fraction__38_comb = {{1{p3_addend_x__11_comb[27]}}, p3_addend_x__11_comb} + {{1{p3_addend_y__11_comb[27]}}, p3_addend_y__11_comb};
  assign p3_abs_fraction__2_comb = p3_fraction__35_comb[28] ? -p3_fraction__35_comb[27:0] : p3_fraction__35_comb[27:0];
  assign p3_abs_fraction__3_comb = p3_fraction__36_comb[28] ? -p3_fraction__36_comb[27:0] : p3_fraction__36_comb[27:0];
  assign p3_abs_fraction__4_comb = p3_fraction__37_comb[28] ? -p3_fraction__37_comb[27:0] : p3_fraction__37_comb[27:0];
  assign p3_abs_fraction__5_comb = p3_fraction__38_comb[28] ? -p3_fraction__38_comb[27:0] : p3_fraction__38_comb[27:0];
  assign p3_reverse_8431_comb = {p3_abs_fraction__2_comb[0], p3_abs_fraction__2_comb[1], p3_abs_fraction__2_comb[2], p3_abs_fraction__2_comb[3], p3_abs_fraction__2_comb[4], p3_abs_fraction__2_comb[5], p3_abs_fraction__2_comb[6], p3_abs_fraction__2_comb[7], p3_abs_fraction__2_comb[8], p3_abs_fraction__2_comb[9], p3_abs_fraction__2_comb[10], p3_abs_fraction__2_comb[11], p3_abs_fraction__2_comb[12], p3_abs_fraction__2_comb[13], p3_abs_fraction__2_comb[14], p3_abs_fraction__2_comb[15], p3_abs_fraction__2_comb[16], p3_abs_fraction__2_comb[17], p3_abs_fraction__2_comb[18], p3_abs_fraction__2_comb[19], p3_abs_fraction__2_comb[20], p3_abs_fraction__2_comb[21], p3_abs_fraction__2_comb[22], p3_abs_fraction__2_comb[23], p3_abs_fraction__2_comb[24], p3_abs_fraction__2_comb[25], p3_abs_fraction__2_comb[26], p3_abs_fraction__2_comb[27]};
  assign p3_reverse_8432_comb = {p3_abs_fraction__3_comb[0], p3_abs_fraction__3_comb[1], p3_abs_fraction__3_comb[2], p3_abs_fraction__3_comb[3], p3_abs_fraction__3_comb[4], p3_abs_fraction__3_comb[5], p3_abs_fraction__3_comb[6], p3_abs_fraction__3_comb[7], p3_abs_fraction__3_comb[8], p3_abs_fraction__3_comb[9], p3_abs_fraction__3_comb[10], p3_abs_fraction__3_comb[11], p3_abs_fraction__3_comb[12], p3_abs_fraction__3_comb[13], p3_abs_fraction__3_comb[14], p3_abs_fraction__3_comb[15], p3_abs_fraction__3_comb[16], p3_abs_fraction__3_comb[17], p3_abs_fraction__3_comb[18], p3_abs_fraction__3_comb[19], p3_abs_fraction__3_comb[20], p3_abs_fraction__3_comb[21], p3_abs_fraction__3_comb[22], p3_abs_fraction__3_comb[23], p3_abs_fraction__3_comb[24], p3_abs_fraction__3_comb[25], p3_abs_fraction__3_comb[26], p3_abs_fraction__3_comb[27]};
  assign p3_reverse_8433_comb = {p3_abs_fraction__4_comb[0], p3_abs_fraction__4_comb[1], p3_abs_fraction__4_comb[2], p3_abs_fraction__4_comb[3], p3_abs_fraction__4_comb[4], p3_abs_fraction__4_comb[5], p3_abs_fraction__4_comb[6], p3_abs_fraction__4_comb[7], p3_abs_fraction__4_comb[8], p3_abs_fraction__4_comb[9], p3_abs_fraction__4_comb[10], p3_abs_fraction__4_comb[11], p3_abs_fraction__4_comb[12], p3_abs_fraction__4_comb[13], p3_abs_fraction__4_comb[14], p3_abs_fraction__4_comb[15], p3_abs_fraction__4_comb[16], p3_abs_fraction__4_comb[17], p3_abs_fraction__4_comb[18], p3_abs_fraction__4_comb[19], p3_abs_fraction__4_comb[20], p3_abs_fraction__4_comb[21], p3_abs_fraction__4_comb[22], p3_abs_fraction__4_comb[23], p3_abs_fraction__4_comb[24], p3_abs_fraction__4_comb[25], p3_abs_fraction__4_comb[26], p3_abs_fraction__4_comb[27]};
  assign p3_reverse_8434_comb = {p3_abs_fraction__5_comb[0], p3_abs_fraction__5_comb[1], p3_abs_fraction__5_comb[2], p3_abs_fraction__5_comb[3], p3_abs_fraction__5_comb[4], p3_abs_fraction__5_comb[5], p3_abs_fraction__5_comb[6], p3_abs_fraction__5_comb[7], p3_abs_fraction__5_comb[8], p3_abs_fraction__5_comb[9], p3_abs_fraction__5_comb[10], p3_abs_fraction__5_comb[11], p3_abs_fraction__5_comb[12], p3_abs_fraction__5_comb[13], p3_abs_fraction__5_comb[14], p3_abs_fraction__5_comb[15], p3_abs_fraction__5_comb[16], p3_abs_fraction__5_comb[17], p3_abs_fraction__5_comb[18], p3_abs_fraction__5_comb[19], p3_abs_fraction__5_comb[20], p3_abs_fraction__5_comb[21], p3_abs_fraction__5_comb[22], p3_abs_fraction__5_comb[23], p3_abs_fraction__5_comb[24], p3_abs_fraction__5_comb[25], p3_abs_fraction__5_comb[26], p3_abs_fraction__5_comb[27]};
  assign p3_one_hot_8435_comb = {p3_reverse_8431_comb[27:0] == 28'h000_0000, p3_reverse_8431_comb[27] && p3_reverse_8431_comb[26:0] == 27'h000_0000, p3_reverse_8431_comb[26] && p3_reverse_8431_comb[25:0] == 26'h000_0000, p3_reverse_8431_comb[25] && p3_reverse_8431_comb[24:0] == 25'h000_0000, p3_reverse_8431_comb[24] && p3_reverse_8431_comb[23:0] == 24'h00_0000, p3_reverse_8431_comb[23] && p3_reverse_8431_comb[22:0] == 23'h00_0000, p3_reverse_8431_comb[22] && p3_reverse_8431_comb[21:0] == 22'h00_0000, p3_reverse_8431_comb[21] && p3_reverse_8431_comb[20:0] == 21'h00_0000, p3_reverse_8431_comb[20] && p3_reverse_8431_comb[19:0] == 20'h0_0000, p3_reverse_8431_comb[19] && p3_reverse_8431_comb[18:0] == 19'h0_0000, p3_reverse_8431_comb[18] && p3_reverse_8431_comb[17:0] == 18'h0_0000, p3_reverse_8431_comb[17] && p3_reverse_8431_comb[16:0] == 17'h0_0000, p3_reverse_8431_comb[16] && p3_reverse_8431_comb[15:0] == 16'h0000, p3_reverse_8431_comb[15] && p3_reverse_8431_comb[14:0] == 15'h0000, p3_reverse_8431_comb[14] && p3_reverse_8431_comb[13:0] == 14'h0000, p3_reverse_8431_comb[13] && p3_reverse_8431_comb[12:0] == 13'h0000, p3_reverse_8431_comb[12] && p3_reverse_8431_comb[11:0] == 12'h000, p3_reverse_8431_comb[11] && p3_reverse_8431_comb[10:0] == 11'h000, p3_reverse_8431_comb[10] && p3_reverse_8431_comb[9:0] == 10'h000, p3_reverse_8431_comb[9] && p3_reverse_8431_comb[8:0] == 9'h000, p3_reverse_8431_comb[8] && p3_reverse_8431_comb[7:0] == 8'h00, p3_reverse_8431_comb[7] && p3_reverse_8431_comb[6:0] == 7'h00, p3_reverse_8431_comb[6] && p3_reverse_8431_comb[5:0] == 6'h00, p3_reverse_8431_comb[5] && p3_reverse_8431_comb[4:0] == 5'h00, p3_reverse_8431_comb[4] && p3_reverse_8431_comb[3:0] == 4'h0, p3_reverse_8431_comb[3] && p3_reverse_8431_comb[2:0] == 3'h0, p3_reverse_8431_comb[2] && p3_reverse_8431_comb[1:0] == 2'h0, p3_reverse_8431_comb[1] && !p3_reverse_8431_comb[0], p3_reverse_8431_comb[0]};
  assign p3_one_hot_8436_comb = {p3_reverse_8432_comb[27:0] == 28'h000_0000, p3_reverse_8432_comb[27] && p3_reverse_8432_comb[26:0] == 27'h000_0000, p3_reverse_8432_comb[26] && p3_reverse_8432_comb[25:0] == 26'h000_0000, p3_reverse_8432_comb[25] && p3_reverse_8432_comb[24:0] == 25'h000_0000, p3_reverse_8432_comb[24] && p3_reverse_8432_comb[23:0] == 24'h00_0000, p3_reverse_8432_comb[23] && p3_reverse_8432_comb[22:0] == 23'h00_0000, p3_reverse_8432_comb[22] && p3_reverse_8432_comb[21:0] == 22'h00_0000, p3_reverse_8432_comb[21] && p3_reverse_8432_comb[20:0] == 21'h00_0000, p3_reverse_8432_comb[20] && p3_reverse_8432_comb[19:0] == 20'h0_0000, p3_reverse_8432_comb[19] && p3_reverse_8432_comb[18:0] == 19'h0_0000, p3_reverse_8432_comb[18] && p3_reverse_8432_comb[17:0] == 18'h0_0000, p3_reverse_8432_comb[17] && p3_reverse_8432_comb[16:0] == 17'h0_0000, p3_reverse_8432_comb[16] && p3_reverse_8432_comb[15:0] == 16'h0000, p3_reverse_8432_comb[15] && p3_reverse_8432_comb[14:0] == 15'h0000, p3_reverse_8432_comb[14] && p3_reverse_8432_comb[13:0] == 14'h0000, p3_reverse_8432_comb[13] && p3_reverse_8432_comb[12:0] == 13'h0000, p3_reverse_8432_comb[12] && p3_reverse_8432_comb[11:0] == 12'h000, p3_reverse_8432_comb[11] && p3_reverse_8432_comb[10:0] == 11'h000, p3_reverse_8432_comb[10] && p3_reverse_8432_comb[9:0] == 10'h000, p3_reverse_8432_comb[9] && p3_reverse_8432_comb[8:0] == 9'h000, p3_reverse_8432_comb[8] && p3_reverse_8432_comb[7:0] == 8'h00, p3_reverse_8432_comb[7] && p3_reverse_8432_comb[6:0] == 7'h00, p3_reverse_8432_comb[6] && p3_reverse_8432_comb[5:0] == 6'h00, p3_reverse_8432_comb[5] && p3_reverse_8432_comb[4:0] == 5'h00, p3_reverse_8432_comb[4] && p3_reverse_8432_comb[3:0] == 4'h0, p3_reverse_8432_comb[3] && p3_reverse_8432_comb[2:0] == 3'h0, p3_reverse_8432_comb[2] && p3_reverse_8432_comb[1:0] == 2'h0, p3_reverse_8432_comb[1] && !p3_reverse_8432_comb[0], p3_reverse_8432_comb[0]};
  assign p3_one_hot_8437_comb = {p3_reverse_8433_comb[27:0] == 28'h000_0000, p3_reverse_8433_comb[27] && p3_reverse_8433_comb[26:0] == 27'h000_0000, p3_reverse_8433_comb[26] && p3_reverse_8433_comb[25:0] == 26'h000_0000, p3_reverse_8433_comb[25] && p3_reverse_8433_comb[24:0] == 25'h000_0000, p3_reverse_8433_comb[24] && p3_reverse_8433_comb[23:0] == 24'h00_0000, p3_reverse_8433_comb[23] && p3_reverse_8433_comb[22:0] == 23'h00_0000, p3_reverse_8433_comb[22] && p3_reverse_8433_comb[21:0] == 22'h00_0000, p3_reverse_8433_comb[21] && p3_reverse_8433_comb[20:0] == 21'h00_0000, p3_reverse_8433_comb[20] && p3_reverse_8433_comb[19:0] == 20'h0_0000, p3_reverse_8433_comb[19] && p3_reverse_8433_comb[18:0] == 19'h0_0000, p3_reverse_8433_comb[18] && p3_reverse_8433_comb[17:0] == 18'h0_0000, p3_reverse_8433_comb[17] && p3_reverse_8433_comb[16:0] == 17'h0_0000, p3_reverse_8433_comb[16] && p3_reverse_8433_comb[15:0] == 16'h0000, p3_reverse_8433_comb[15] && p3_reverse_8433_comb[14:0] == 15'h0000, p3_reverse_8433_comb[14] && p3_reverse_8433_comb[13:0] == 14'h0000, p3_reverse_8433_comb[13] && p3_reverse_8433_comb[12:0] == 13'h0000, p3_reverse_8433_comb[12] && p3_reverse_8433_comb[11:0] == 12'h000, p3_reverse_8433_comb[11] && p3_reverse_8433_comb[10:0] == 11'h000, p3_reverse_8433_comb[10] && p3_reverse_8433_comb[9:0] == 10'h000, p3_reverse_8433_comb[9] && p3_reverse_8433_comb[8:0] == 9'h000, p3_reverse_8433_comb[8] && p3_reverse_8433_comb[7:0] == 8'h00, p3_reverse_8433_comb[7] && p3_reverse_8433_comb[6:0] == 7'h00, p3_reverse_8433_comb[6] && p3_reverse_8433_comb[5:0] == 6'h00, p3_reverse_8433_comb[5] && p3_reverse_8433_comb[4:0] == 5'h00, p3_reverse_8433_comb[4] && p3_reverse_8433_comb[3:0] == 4'h0, p3_reverse_8433_comb[3] && p3_reverse_8433_comb[2:0] == 3'h0, p3_reverse_8433_comb[2] && p3_reverse_8433_comb[1:0] == 2'h0, p3_reverse_8433_comb[1] && !p3_reverse_8433_comb[0], p3_reverse_8433_comb[0]};
  assign p3_one_hot_8438_comb = {p3_reverse_8434_comb[27:0] == 28'h000_0000, p3_reverse_8434_comb[27] && p3_reverse_8434_comb[26:0] == 27'h000_0000, p3_reverse_8434_comb[26] && p3_reverse_8434_comb[25:0] == 26'h000_0000, p3_reverse_8434_comb[25] && p3_reverse_8434_comb[24:0] == 25'h000_0000, p3_reverse_8434_comb[24] && p3_reverse_8434_comb[23:0] == 24'h00_0000, p3_reverse_8434_comb[23] && p3_reverse_8434_comb[22:0] == 23'h00_0000, p3_reverse_8434_comb[22] && p3_reverse_8434_comb[21:0] == 22'h00_0000, p3_reverse_8434_comb[21] && p3_reverse_8434_comb[20:0] == 21'h00_0000, p3_reverse_8434_comb[20] && p3_reverse_8434_comb[19:0] == 20'h0_0000, p3_reverse_8434_comb[19] && p3_reverse_8434_comb[18:0] == 19'h0_0000, p3_reverse_8434_comb[18] && p3_reverse_8434_comb[17:0] == 18'h0_0000, p3_reverse_8434_comb[17] && p3_reverse_8434_comb[16:0] == 17'h0_0000, p3_reverse_8434_comb[16] && p3_reverse_8434_comb[15:0] == 16'h0000, p3_reverse_8434_comb[15] && p3_reverse_8434_comb[14:0] == 15'h0000, p3_reverse_8434_comb[14] && p3_reverse_8434_comb[13:0] == 14'h0000, p3_reverse_8434_comb[13] && p3_reverse_8434_comb[12:0] == 13'h0000, p3_reverse_8434_comb[12] && p3_reverse_8434_comb[11:0] == 12'h000, p3_reverse_8434_comb[11] && p3_reverse_8434_comb[10:0] == 11'h000, p3_reverse_8434_comb[10] && p3_reverse_8434_comb[9:0] == 10'h000, p3_reverse_8434_comb[9] && p3_reverse_8434_comb[8:0] == 9'h000, p3_reverse_8434_comb[8] && p3_reverse_8434_comb[7:0] == 8'h00, p3_reverse_8434_comb[7] && p3_reverse_8434_comb[6:0] == 7'h00, p3_reverse_8434_comb[6] && p3_reverse_8434_comb[5:0] == 6'h00, p3_reverse_8434_comb[5] && p3_reverse_8434_comb[4:0] == 5'h00, p3_reverse_8434_comb[4] && p3_reverse_8434_comb[3:0] == 4'h0, p3_reverse_8434_comb[3] && p3_reverse_8434_comb[2:0] == 3'h0, p3_reverse_8434_comb[2] && p3_reverse_8434_comb[1:0] == 2'h0, p3_reverse_8434_comb[1] && !p3_reverse_8434_comb[0], p3_reverse_8434_comb[0]};
  assign p3_encode_8439_comb = {p3_one_hot_8435_comb[16] | p3_one_hot_8435_comb[17] | p3_one_hot_8435_comb[18] | p3_one_hot_8435_comb[19] | p3_one_hot_8435_comb[20] | p3_one_hot_8435_comb[21] | p3_one_hot_8435_comb[22] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[24] | p3_one_hot_8435_comb[25] | p3_one_hot_8435_comb[26] | p3_one_hot_8435_comb[27] | p3_one_hot_8435_comb[28], p3_one_hot_8435_comb[8] | p3_one_hot_8435_comb[9] | p3_one_hot_8435_comb[10] | p3_one_hot_8435_comb[11] | p3_one_hot_8435_comb[12] | p3_one_hot_8435_comb[13] | p3_one_hot_8435_comb[14] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[24] | p3_one_hot_8435_comb[25] | p3_one_hot_8435_comb[26] | p3_one_hot_8435_comb[27] | p3_one_hot_8435_comb[28], p3_one_hot_8435_comb[4] | p3_one_hot_8435_comb[5] | p3_one_hot_8435_comb[6] | p3_one_hot_8435_comb[7] | p3_one_hot_8435_comb[12] | p3_one_hot_8435_comb[13] | p3_one_hot_8435_comb[14] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[20] | p3_one_hot_8435_comb[21] | p3_one_hot_8435_comb[22] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[28], p3_one_hot_8435_comb[2] | p3_one_hot_8435_comb[3] | p3_one_hot_8435_comb[6] | p3_one_hot_8435_comb[7] | p3_one_hot_8435_comb[10] | p3_one_hot_8435_comb[11] | p3_one_hot_8435_comb[14] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[18] | p3_one_hot_8435_comb[19] | p3_one_hot_8435_comb[22] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[26] | p3_one_hot_8435_comb[27], p3_one_hot_8435_comb[1] | p3_one_hot_8435_comb[3] | p3_one_hot_8435_comb[5] | p3_one_hot_8435_comb[7] | p3_one_hot_8435_comb[9] | p3_one_hot_8435_comb[11] | p3_one_hot_8435_comb[13] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[17] | p3_one_hot_8435_comb[19] | p3_one_hot_8435_comb[21] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[25] | p3_one_hot_8435_comb[27]};
  assign p3_encode_8440_comb = {p3_one_hot_8436_comb[16] | p3_one_hot_8436_comb[17] | p3_one_hot_8436_comb[18] | p3_one_hot_8436_comb[19] | p3_one_hot_8436_comb[20] | p3_one_hot_8436_comb[21] | p3_one_hot_8436_comb[22] | p3_one_hot_8436_comb[23] | p3_one_hot_8436_comb[24] | p3_one_hot_8436_comb[25] | p3_one_hot_8436_comb[26] | p3_one_hot_8436_comb[27] | p3_one_hot_8436_comb[28], p3_one_hot_8436_comb[8] | p3_one_hot_8436_comb[9] | p3_one_hot_8436_comb[10] | p3_one_hot_8436_comb[11] | p3_one_hot_8436_comb[12] | p3_one_hot_8436_comb[13] | p3_one_hot_8436_comb[14] | p3_one_hot_8436_comb[15] | p3_one_hot_8436_comb[24] | p3_one_hot_8436_comb[25] | p3_one_hot_8436_comb[26] | p3_one_hot_8436_comb[27] | p3_one_hot_8436_comb[28], p3_one_hot_8436_comb[4] | p3_one_hot_8436_comb[5] | p3_one_hot_8436_comb[6] | p3_one_hot_8436_comb[7] | p3_one_hot_8436_comb[12] | p3_one_hot_8436_comb[13] | p3_one_hot_8436_comb[14] | p3_one_hot_8436_comb[15] | p3_one_hot_8436_comb[20] | p3_one_hot_8436_comb[21] | p3_one_hot_8436_comb[22] | p3_one_hot_8436_comb[23] | p3_one_hot_8436_comb[28], p3_one_hot_8436_comb[2] | p3_one_hot_8436_comb[3] | p3_one_hot_8436_comb[6] | p3_one_hot_8436_comb[7] | p3_one_hot_8436_comb[10] | p3_one_hot_8436_comb[11] | p3_one_hot_8436_comb[14] | p3_one_hot_8436_comb[15] | p3_one_hot_8436_comb[18] | p3_one_hot_8436_comb[19] | p3_one_hot_8436_comb[22] | p3_one_hot_8436_comb[23] | p3_one_hot_8436_comb[26] | p3_one_hot_8436_comb[27], p3_one_hot_8436_comb[1] | p3_one_hot_8436_comb[3] | p3_one_hot_8436_comb[5] | p3_one_hot_8436_comb[7] | p3_one_hot_8436_comb[9] | p3_one_hot_8436_comb[11] | p3_one_hot_8436_comb[13] | p3_one_hot_8436_comb[15] | p3_one_hot_8436_comb[17] | p3_one_hot_8436_comb[19] | p3_one_hot_8436_comb[21] | p3_one_hot_8436_comb[23] | p3_one_hot_8436_comb[25] | p3_one_hot_8436_comb[27]};
  assign p3_encode_8441_comb = {p3_one_hot_8437_comb[16] | p3_one_hot_8437_comb[17] | p3_one_hot_8437_comb[18] | p3_one_hot_8437_comb[19] | p3_one_hot_8437_comb[20] | p3_one_hot_8437_comb[21] | p3_one_hot_8437_comb[22] | p3_one_hot_8437_comb[23] | p3_one_hot_8437_comb[24] | p3_one_hot_8437_comb[25] | p3_one_hot_8437_comb[26] | p3_one_hot_8437_comb[27] | p3_one_hot_8437_comb[28], p3_one_hot_8437_comb[8] | p3_one_hot_8437_comb[9] | p3_one_hot_8437_comb[10] | p3_one_hot_8437_comb[11] | p3_one_hot_8437_comb[12] | p3_one_hot_8437_comb[13] | p3_one_hot_8437_comb[14] | p3_one_hot_8437_comb[15] | p3_one_hot_8437_comb[24] | p3_one_hot_8437_comb[25] | p3_one_hot_8437_comb[26] | p3_one_hot_8437_comb[27] | p3_one_hot_8437_comb[28], p3_one_hot_8437_comb[4] | p3_one_hot_8437_comb[5] | p3_one_hot_8437_comb[6] | p3_one_hot_8437_comb[7] | p3_one_hot_8437_comb[12] | p3_one_hot_8437_comb[13] | p3_one_hot_8437_comb[14] | p3_one_hot_8437_comb[15] | p3_one_hot_8437_comb[20] | p3_one_hot_8437_comb[21] | p3_one_hot_8437_comb[22] | p3_one_hot_8437_comb[23] | p3_one_hot_8437_comb[28], p3_one_hot_8437_comb[2] | p3_one_hot_8437_comb[3] | p3_one_hot_8437_comb[6] | p3_one_hot_8437_comb[7] | p3_one_hot_8437_comb[10] | p3_one_hot_8437_comb[11] | p3_one_hot_8437_comb[14] | p3_one_hot_8437_comb[15] | p3_one_hot_8437_comb[18] | p3_one_hot_8437_comb[19] | p3_one_hot_8437_comb[22] | p3_one_hot_8437_comb[23] | p3_one_hot_8437_comb[26] | p3_one_hot_8437_comb[27], p3_one_hot_8437_comb[1] | p3_one_hot_8437_comb[3] | p3_one_hot_8437_comb[5] | p3_one_hot_8437_comb[7] | p3_one_hot_8437_comb[9] | p3_one_hot_8437_comb[11] | p3_one_hot_8437_comb[13] | p3_one_hot_8437_comb[15] | p3_one_hot_8437_comb[17] | p3_one_hot_8437_comb[19] | p3_one_hot_8437_comb[21] | p3_one_hot_8437_comb[23] | p3_one_hot_8437_comb[25] | p3_one_hot_8437_comb[27]};
  assign p3_encode_8442_comb = {p3_one_hot_8438_comb[16] | p3_one_hot_8438_comb[17] | p3_one_hot_8438_comb[18] | p3_one_hot_8438_comb[19] | p3_one_hot_8438_comb[20] | p3_one_hot_8438_comb[21] | p3_one_hot_8438_comb[22] | p3_one_hot_8438_comb[23] | p3_one_hot_8438_comb[24] | p3_one_hot_8438_comb[25] | p3_one_hot_8438_comb[26] | p3_one_hot_8438_comb[27] | p3_one_hot_8438_comb[28], p3_one_hot_8438_comb[8] | p3_one_hot_8438_comb[9] | p3_one_hot_8438_comb[10] | p3_one_hot_8438_comb[11] | p3_one_hot_8438_comb[12] | p3_one_hot_8438_comb[13] | p3_one_hot_8438_comb[14] | p3_one_hot_8438_comb[15] | p3_one_hot_8438_comb[24] | p3_one_hot_8438_comb[25] | p3_one_hot_8438_comb[26] | p3_one_hot_8438_comb[27] | p3_one_hot_8438_comb[28], p3_one_hot_8438_comb[4] | p3_one_hot_8438_comb[5] | p3_one_hot_8438_comb[6] | p3_one_hot_8438_comb[7] | p3_one_hot_8438_comb[12] | p3_one_hot_8438_comb[13] | p3_one_hot_8438_comb[14] | p3_one_hot_8438_comb[15] | p3_one_hot_8438_comb[20] | p3_one_hot_8438_comb[21] | p3_one_hot_8438_comb[22] | p3_one_hot_8438_comb[23] | p3_one_hot_8438_comb[28], p3_one_hot_8438_comb[2] | p3_one_hot_8438_comb[3] | p3_one_hot_8438_comb[6] | p3_one_hot_8438_comb[7] | p3_one_hot_8438_comb[10] | p3_one_hot_8438_comb[11] | p3_one_hot_8438_comb[14] | p3_one_hot_8438_comb[15] | p3_one_hot_8438_comb[18] | p3_one_hot_8438_comb[19] | p3_one_hot_8438_comb[22] | p3_one_hot_8438_comb[23] | p3_one_hot_8438_comb[26] | p3_one_hot_8438_comb[27], p3_one_hot_8438_comb[1] | p3_one_hot_8438_comb[3] | p3_one_hot_8438_comb[5] | p3_one_hot_8438_comb[7] | p3_one_hot_8438_comb[9] | p3_one_hot_8438_comb[11] | p3_one_hot_8438_comb[13] | p3_one_hot_8438_comb[15] | p3_one_hot_8438_comb[17] | p3_one_hot_8438_comb[19] | p3_one_hot_8438_comb[21] | p3_one_hot_8438_comb[23] | p3_one_hot_8438_comb[25] | p3_one_hot_8438_comb[27]};
  assign p3_carry_bit__2_comb = p3_abs_fraction__2_comb[27];
  assign p3_cancel__2_comb = p3_encode_8439_comb[1] | p3_encode_8439_comb[2] | p3_encode_8439_comb[3] | p3_encode_8439_comb[4];
  assign p3_carry_bit__3_comb = p3_abs_fraction__3_comb[27];
  assign p3_cancel__3_comb = p3_encode_8440_comb[1] | p3_encode_8440_comb[2] | p3_encode_8440_comb[3] | p3_encode_8440_comb[4];
  assign p3_carry_bit__4_comb = p3_abs_fraction__4_comb[27];
  assign p3_cancel__4_comb = p3_encode_8441_comb[1] | p3_encode_8441_comb[2] | p3_encode_8441_comb[3] | p3_encode_8441_comb[4];
  assign p3_carry_bit__5_comb = p3_abs_fraction__5_comb[27];
  assign p3_cancel__5_comb = p3_encode_8442_comb[1] | p3_encode_8442_comb[2] | p3_encode_8442_comb[3] | p3_encode_8442_comb[4];
  assign p3_leading_zeroes__2_comb = {23'h00_0000, p3_encode_8439_comb};
  assign p3_leading_zeroes__3_comb = {23'h00_0000, p3_encode_8440_comb};
  assign p3_leading_zeroes__4_comb = {23'h00_0000, p3_encode_8441_comb};
  assign p3_leading_zeroes__5_comb = {23'h00_0000, p3_encode_8442_comb};
  assign p3_and_8495_comb = ~p3_carry_bit__2_comb & ~p3_cancel__2_comb;
  assign p3_and_8496_comb = ~p3_carry_bit__2_comb & p3_cancel__2_comb;
  assign p3_and_8497_comb = p3_carry_bit__2_comb & ~p3_cancel__2_comb;
  assign p3_carry_fraction__4_comb = p3_abs_fraction__2_comb[27:1];
  assign p3_add_8501_comb = p3_leading_zeroes__2_comb + 28'hfff_ffff;
  assign p3_and_8502_comb = ~p3_carry_bit__3_comb & ~p3_cancel__3_comb;
  assign p3_and_8503_comb = ~p3_carry_bit__3_comb & p3_cancel__3_comb;
  assign p3_and_8504_comb = p3_carry_bit__3_comb & ~p3_cancel__3_comb;
  assign p3_carry_fraction__6_comb = p3_abs_fraction__3_comb[27:1];
  assign p3_add_8508_comb = p3_leading_zeroes__3_comb + 28'hfff_ffff;
  assign p3_and_8509_comb = ~p3_carry_bit__4_comb & ~p3_cancel__4_comb;
  assign p3_and_8510_comb = ~p3_carry_bit__4_comb & p3_cancel__4_comb;
  assign p3_and_8511_comb = p3_carry_bit__4_comb & ~p3_cancel__4_comb;
  assign p3_carry_fraction__8_comb = p3_abs_fraction__4_comb[27:1];
  assign p3_add_8515_comb = p3_leading_zeroes__4_comb + 28'hfff_ffff;
  assign p3_and_8516_comb = ~p3_carry_bit__5_comb & ~p3_cancel__5_comb;
  assign p3_and_8517_comb = ~p3_carry_bit__5_comb & p3_cancel__5_comb;
  assign p3_and_8518_comb = p3_carry_bit__5_comb & ~p3_cancel__5_comb;
  assign p3_carry_fraction__10_comb = p3_abs_fraction__5_comb[27:1];
  assign p3_add_8522_comb = p3_leading_zeroes__5_comb + 28'hfff_ffff;
  assign p3_concat_8523_comb = {p3_and_8495_comb, p3_and_8496_comb, p3_and_8497_comb};
  assign p3_carry_fraction__5_comb = p3_carry_fraction__4_comb | {26'h000_0000, p3_abs_fraction__2_comb[0]};
  assign p3_cancel_fraction__2_comb = p3_add_8501_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__2_comb[26:0] << p3_add_8501_comb;
  assign p3_concat_8526_comb = {p3_and_8502_comb, p3_and_8503_comb, p3_and_8504_comb};
  assign p3_carry_fraction__7_comb = p3_carry_fraction__6_comb | {26'h000_0000, p3_abs_fraction__3_comb[0]};
  assign p3_cancel_fraction__3_comb = p3_add_8508_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__3_comb[26:0] << p3_add_8508_comb;
  assign p3_concat_8529_comb = {p3_and_8509_comb, p3_and_8510_comb, p3_and_8511_comb};
  assign p3_carry_fraction__9_comb = p3_carry_fraction__8_comb | {26'h000_0000, p3_abs_fraction__4_comb[0]};
  assign p3_cancel_fraction__4_comb = p3_add_8515_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__4_comb[26:0] << p3_add_8515_comb;
  assign p3_concat_8532_comb = {p3_and_8516_comb, p3_and_8517_comb, p3_and_8518_comb};
  assign p3_carry_fraction__11_comb = p3_carry_fraction__10_comb | {26'h000_0000, p3_abs_fraction__5_comb[0]};
  assign p3_cancel_fraction__5_comb = p3_add_8522_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__5_comb[26:0] << p3_add_8522_comb;
  assign p3_shifted_fraction__2_comb = p3_carry_fraction__5_comb & {27{p3_concat_8523_comb[0]}} | p3_cancel_fraction__2_comb & {27{p3_concat_8523_comb[1]}} | p3_abs_fraction__2_comb[26:0] & {27{p3_concat_8523_comb[2]}};
  assign p3_shifted_fraction__3_comb = p3_carry_fraction__7_comb & {27{p3_concat_8526_comb[0]}} | p3_cancel_fraction__3_comb & {27{p3_concat_8526_comb[1]}} | p3_abs_fraction__3_comb[26:0] & {27{p3_concat_8526_comb[2]}};
  assign p3_shifted_fraction__4_comb = p3_carry_fraction__9_comb & {27{p3_concat_8529_comb[0]}} | p3_cancel_fraction__4_comb & {27{p3_concat_8529_comb[1]}} | p3_abs_fraction__4_comb[26:0] & {27{p3_concat_8529_comb[2]}};
  assign p3_shifted_fraction__5_comb = p3_carry_fraction__11_comb & {27{p3_concat_8532_comb[0]}} | p3_cancel_fraction__5_comb & {27{p3_concat_8532_comb[1]}} | p3_abs_fraction__5_comb[26:0] & {27{p3_concat_8532_comb[2]}};
  assign p3_normal_chunk__2_comb = p3_shifted_fraction__2_comb[2:0];
  assign p3_half_way_chunk__2_comb = p3_shifted_fraction__2_comb[3:2];
  assign p3_normal_chunk__3_comb = p3_shifted_fraction__3_comb[2:0];
  assign p3_half_way_chunk__3_comb = p3_shifted_fraction__3_comb[3:2];
  assign p3_normal_chunk__4_comb = p3_shifted_fraction__4_comb[2:0];
  assign p3_half_way_chunk__4_comb = p3_shifted_fraction__4_comb[3:2];
  assign p3_normal_chunk__5_comb = p3_shifted_fraction__5_comb[2:0];
  assign p3_half_way_chunk__5_comb = p3_shifted_fraction__5_comb[3:2];
  assign p3_add_8574_comb = {1'h0, p3_shifted_fraction__2_comb[26:3]} + 25'h000_0001;
  assign p3_add_8578_comb = {1'h0, p3_shifted_fraction__3_comb[26:3]} + 25'h000_0001;
  assign p3_add_8582_comb = {1'h0, p3_shifted_fraction__4_comb[26:3]} + 25'h000_0001;
  assign p3_add_8586_comb = {1'h0, p3_shifted_fraction__5_comb[26:3]} + 25'h000_0001;
  assign p3_do_round_up__7_comb = p3_normal_chunk__2_comb > 3'h4 | p3_half_way_chunk__2_comb == 2'h3;
  assign p3_do_round_up__8_comb = p3_normal_chunk__3_comb > 3'h4 | p3_half_way_chunk__3_comb == 2'h3;
  assign p3_do_round_up__9_comb = p3_normal_chunk__4_comb > 3'h4 | p3_half_way_chunk__4_comb == 2'h3;
  assign p3_do_round_up__10_comb = p3_normal_chunk__5_comb > 3'h4 | p3_half_way_chunk__5_comb == 2'h3;
  assign p3_rounded_fraction__2_comb = p3_do_round_up__7_comb ? {p3_add_8574_comb, p3_normal_chunk__2_comb} : {1'h0, p3_shifted_fraction__2_comb};
  assign p3_rounded_fraction__3_comb = p3_do_round_up__8_comb ? {p3_add_8578_comb, p3_normal_chunk__3_comb} : {1'h0, p3_shifted_fraction__3_comb};
  assign p3_rounded_fraction__4_comb = p3_do_round_up__9_comb ? {p3_add_8582_comb, p3_normal_chunk__4_comb} : {1'h0, p3_shifted_fraction__4_comb};
  assign p3_rounded_fraction__5_comb = p3_do_round_up__10_comb ? {p3_add_8586_comb, p3_normal_chunk__5_comb} : {1'h0, p3_shifted_fraction__5_comb};
  assign p3_rounding_carry__2_comb = p3_rounded_fraction__2_comb[27];
  assign p3_rounding_carry__3_comb = p3_rounded_fraction__3_comb[27];
  assign p3_rounding_carry__4_comb = p3_rounded_fraction__4_comb[27];
  assign p3_rounding_carry__5_comb = p3_rounded_fraction__5_comb[27];
  assign p3_concat_8613_comb = {1'h0, p2_greater_exp_bexp__2};
  assign p3_concat_8615_comb = {1'h0, p2_greater_exp_bexp__3};
  assign p3_add_8620_comb = p3_concat_8613_comb + {8'h00, p3_rounding_carry__2_comb};
  assign p3_add_8622_comb = p3_concat_8615_comb + {8'h00, p3_rounding_carry__3_comb};
  assign p3_add_8624_comb = p3_concat_8613_comb + {8'h00, p3_rounding_carry__4_comb};
  assign p3_add_8626_comb = p3_concat_8615_comb + {8'h00, p3_rounding_carry__5_comb};
  assign p3_add_8643_comb = {1'h0, p3_add_8620_comb} + 10'h001;
  assign p3_add_8646_comb = {1'h0, p3_add_8622_comb} + 10'h001;
  assign p3_add_8649_comb = {1'h0, p3_add_8624_comb} + 10'h001;
  assign p3_add_8652_comb = {1'h0, p3_add_8626_comb} + 10'h001;
  assign p3_wide_exponent__6_comb = p3_add_8643_comb - {5'h00, p3_encode_8439_comb};
  assign p3_wide_exponent__9_comb = p3_add_8646_comb - {5'h00, p3_encode_8440_comb};
  assign p3_wide_exponent__12_comb = p3_add_8649_comb - {5'h00, p3_encode_8441_comb};
  assign p3_wide_exponent__15_comb = p3_add_8652_comb - {5'h00, p3_encode_8442_comb};
  assign p3_wide_exponent__7_comb = p3_wide_exponent__6_comb & {10{p3_fraction__35_comb != 29'h0000_0000}};
  assign p3_wide_exponent__10_comb = p3_wide_exponent__9_comb & {10{p3_fraction__36_comb != 29'h0000_0000}};
  assign p3_wide_exponent__13_comb = p3_wide_exponent__12_comb & {10{p3_fraction__37_comb != 29'h0000_0000}};
  assign p3_wide_exponent__16_comb = p3_wide_exponent__15_comb & {10{p3_fraction__38_comb != 29'h0000_0000}};
  assign p3_wide_exponent__8_comb = p3_wide_exponent__7_comb[8:0] & {9{~p3_wide_exponent__7_comb[9]}};
  assign p3_wide_exponent__11_comb = p3_wide_exponent__10_comb[8:0] & {9{~p3_wide_exponent__10_comb[9]}};
  assign p3_wide_exponent__14_comb = p3_wide_exponent__13_comb[8:0] & {9{~p3_wide_exponent__13_comb[9]}};
  assign p3_wide_exponent__17_comb = p3_wide_exponent__16_comb[8:0] & {9{~p3_wide_exponent__16_comb[9]}};
  assign p3_fraction_is_zero__2_comb = p3_fraction__35_comb == 29'h0000_0000;
  assign p3_add_8747_comb = {2'h0, p3_rounding_carry__2_comb} + 3'h3;
  assign p3_fraction_is_zero__3_comb = p3_fraction__36_comb == 29'h0000_0000;
  assign p3_add_8753_comb = {2'h0, p3_rounding_carry__3_comb} + 3'h3;
  assign p3_fraction_is_zero__4_comb = p3_fraction__37_comb == 29'h0000_0000;
  assign p3_add_8759_comb = {2'h0, p3_rounding_carry__4_comb} + 3'h3;
  assign p3_fraction_is_zero__5_comb = p3_fraction__38_comb == 29'h0000_0000;
  assign p3_add_8765_comb = {2'h0, p3_rounding_carry__5_comb} + 3'h3;
  assign p3_nor_8769_comb = ~(p3_wide_exponent__8_comb[8] | p3_wide_exponent__8_comb[0] & p3_wide_exponent__8_comb[1] & p3_wide_exponent__8_comb[2] & p3_wide_exponent__8_comb[3] & p3_wide_exponent__8_comb[4] & p3_wide_exponent__8_comb[5] & p3_wide_exponent__8_comb[6] & p3_wide_exponent__8_comb[7]);
  assign p3_shrl_8770_comb = p3_rounded_fraction__2_comb >> p3_add_8747_comb;
  assign p3_nor_8774_comb = ~(p3_wide_exponent__11_comb[8] | p3_wide_exponent__11_comb[0] & p3_wide_exponent__11_comb[1] & p3_wide_exponent__11_comb[2] & p3_wide_exponent__11_comb[3] & p3_wide_exponent__11_comb[4] & p3_wide_exponent__11_comb[5] & p3_wide_exponent__11_comb[6] & p3_wide_exponent__11_comb[7]);
  assign p3_shrl_8775_comb = p3_rounded_fraction__3_comb >> p3_add_8753_comb;
  assign p3_nor_8779_comb = ~(p3_wide_exponent__14_comb[8] | p3_wide_exponent__14_comb[0] & p3_wide_exponent__14_comb[1] & p3_wide_exponent__14_comb[2] & p3_wide_exponent__14_comb[3] & p3_wide_exponent__14_comb[4] & p3_wide_exponent__14_comb[5] & p3_wide_exponent__14_comb[6] & p3_wide_exponent__14_comb[7]);
  assign p3_shrl_8780_comb = p3_rounded_fraction__4_comb >> p3_add_8759_comb;
  assign p3_nor_8784_comb = ~(p3_wide_exponent__17_comb[8] | p3_wide_exponent__17_comb[0] & p3_wide_exponent__17_comb[1] & p3_wide_exponent__17_comb[2] & p3_wide_exponent__17_comb[3] & p3_wide_exponent__17_comb[4] & p3_wide_exponent__17_comb[5] & p3_wide_exponent__17_comb[6] & p3_wide_exponent__17_comb[7]);
  assign p3_shrl_8785_comb = p3_rounded_fraction__5_comb >> p3_add_8765_comb;
  assign p3_result_sign__15_comb = ~(~p3_fraction__35_comb[28] | p3_greater_exp_sign__2_comb) | ~(p3_fraction__35_comb[28] | p3_fraction_is_zero__2_comb | ~p3_greater_exp_sign__2_comb);
  assign p3_result_fraction__19_comb = p3_shrl_8770_comb[22:0];
  assign p3_sign_ext_8792_comb = {23{p2_nor_8298}};
  assign p3_result_sign__17_comb = ~(~p3_fraction__36_comb[28] | p3_greater_exp_sign__3_comb) | ~(p3_fraction__36_comb[28] | p3_fraction_is_zero__3_comb | ~p3_greater_exp_sign__3_comb);
  assign p3_result_fraction__21_comb = p3_shrl_8775_comb[22:0];
  assign p3_sign_ext_8798_comb = {23{p2_nor_8302}};
  assign p3_result_sign__20_comb = ~(~p3_fraction__37_comb[28] | p3_greater_exp_sign__4_comb) | ~(p3_fraction__37_comb[28] | p3_fraction_is_zero__4_comb | ~p3_greater_exp_sign__4_comb);
  assign p3_result_fraction__24_comb = p3_shrl_8780_comb[22:0];
  assign p3_result_sign__23_comb = ~(~p3_fraction__38_comb[28] | p3_greater_exp_sign__5_comb) | ~(p3_fraction__38_comb[28] | p3_fraction_is_zero__5_comb | ~p3_greater_exp_sign__5_comb);
  assign p3_result_fraction__27_comb = p3_shrl_8785_comb[22:0];
  assign p3_result_sign__16_comb = p2_is_operand_inf__2 ? p2_not_8307 : p3_result_sign__15_comb;
  assign p3_high_exp__42_comb = 8'hff;
  assign p3_result_fraction__20_comb = p3_result_fraction__19_comb & {23{~(~(p3_wide_exponent__8_comb[1] | p3_wide_exponent__8_comb[2] | p3_wide_exponent__8_comb[3] | p3_wide_exponent__8_comb[4] | p3_wide_exponent__8_comb[5] | p3_wide_exponent__8_comb[6] | p3_wide_exponent__8_comb[7] | p3_wide_exponent__8_comb[8] | p3_wide_exponent__8_comb[0]))}} & {23{p3_nor_8769_comb}} & p3_sign_ext_8792_comb;
  assign p3_nan_fraction__16_comb = 23'h40_0000;
  assign p3_result_sign__18_comb = p2_is_operand_inf__3 ? p2_not_8310 : p3_result_sign__17_comb;
  assign p3_high_exp__43_comb = 8'hff;
  assign p3_result_fraction__22_comb = p3_result_fraction__21_comb & {23{~(~(p3_wide_exponent__11_comb[1] | p3_wide_exponent__11_comb[2] | p3_wide_exponent__11_comb[3] | p3_wide_exponent__11_comb[4] | p3_wide_exponent__11_comb[5] | p3_wide_exponent__11_comb[6] | p3_wide_exponent__11_comb[7] | p3_wide_exponent__11_comb[8] | p3_wide_exponent__11_comb[0]))}} & {23{p3_nor_8774_comb}} & p3_sign_ext_8798_comb;
  assign p3_nan_fraction__17_comb = 23'h40_0000;
  assign p3_result_sign__21_comb = p2_is_operand_inf__2 ? p2_not_8312 : p3_result_sign__20_comb;
  assign p3_high_exp__44_comb = 8'hff;
  assign p3_result_fraction__25_comb = p3_result_fraction__24_comb & {23{~(~(p3_wide_exponent__14_comb[1] | p3_wide_exponent__14_comb[2] | p3_wide_exponent__14_comb[3] | p3_wide_exponent__14_comb[4] | p3_wide_exponent__14_comb[5] | p3_wide_exponent__14_comb[6] | p3_wide_exponent__14_comb[7] | p3_wide_exponent__14_comb[8] | p3_wide_exponent__14_comb[0]))}} & {23{p3_nor_8779_comb}} & p3_sign_ext_8792_comb;
  assign p3_nan_fraction__18_comb = 23'h40_0000;
  assign p3_result_sign__24_comb = p2_is_operand_inf__3 ? p2_not_8314 : p3_result_sign__23_comb;
  assign p3_high_exp__45_comb = 8'hff;
  assign p3_result_fraction__28_comb = p3_result_fraction__27_comb & {23{~(~(p3_wide_exponent__17_comb[1] | p3_wide_exponent__17_comb[2] | p3_wide_exponent__17_comb[3] | p3_wide_exponent__17_comb[4] | p3_wide_exponent__17_comb[5] | p3_wide_exponent__17_comb[6] | p3_wide_exponent__17_comb[7] | p3_wide_exponent__17_comb[8] | p3_wide_exponent__17_comb[0]))}} & {23{p3_nor_8784_comb}} & p3_sign_ext_8798_comb;
  assign p3_nan_fraction__19_comb = 23'h40_0000;
  assign p3_result_sign__19_comb = ~p2_is_result_nan__7 & p3_result_sign__16_comb;
  assign p3_result_exponent__3_comb = p2_is_result_nan__7 | p2_is_operand_inf__2 | ~p3_nor_8769_comb ? p3_high_exp__42_comb : p3_wide_exponent__8_comb[7:0];
  assign p3_result_fraction__23_comb = p2_is_result_nan__7 ? p3_nan_fraction__16_comb : p3_result_fraction__20_comb;
  assign p3_result_sign__22_comb = ~p2_is_result_nan__8 & p3_result_sign__18_comb;
  assign p3_result_exponent__4_comb = p2_is_result_nan__8 | p2_is_operand_inf__3 | ~p3_nor_8774_comb ? p3_high_exp__43_comb : p3_wide_exponent__11_comb[7:0];
  assign p3_result_fraction__26_comb = p2_is_result_nan__8 ? p3_nan_fraction__17_comb : p3_result_fraction__22_comb;
  assign p3_result_sign__25_comb = ~p2_is_result_nan__9 & p3_result_sign__21_comb;
  assign p3_result_exponent__5_comb = p2_is_result_nan__9 | p2_is_operand_inf__2 | ~p3_nor_8779_comb ? p3_high_exp__44_comb : p3_wide_exponent__14_comb[7:0];
  assign p3_result_fraction__29_comb = p2_is_result_nan__9 ? p3_nan_fraction__18_comb : p3_result_fraction__25_comb;
  assign p3_result_sign__26_comb = ~p2_is_result_nan__10 & p3_result_sign__24_comb;
  assign p3_result_exponent__6_comb = p2_is_result_nan__10 | p2_is_operand_inf__3 | ~p3_nor_8784_comb ? p3_high_exp__45_comb : p3_wide_exponent__17_comb[7:0];
  assign p3_result_fraction__30_comb = p2_is_result_nan__10 ? p3_nan_fraction__19_comb : p3_result_fraction__28_comb;
  assign p3_out0_r_comb = {p3_result_sign__19_comb, p3_result_exponent__3_comb, p3_result_fraction__23_comb};
  assign p3_out0_i_comb = {p3_result_sign__22_comb, p3_result_exponent__4_comb, p3_result_fraction__26_comb};
  assign p3_out1_r_comb = {p3_result_sign__25_comb, p3_result_exponent__5_comb, p3_result_fraction__29_comb};
  assign p3_out1_i_comb = {p3_result_sign__26_comb, p3_result_exponent__6_comb, p3_result_fraction__30_comb};
  assign p3_tuple_8861_comb = {p3_out0_r_comb, p3_out0_i_comb, p3_out1_r_comb, p3_out1_i_comb};

  // Registers for pipe stage 3:
  reg [127:0] p3_tuple_8861;
  always_ff @ (posedge clk) begin
    p3_tuple_8861 <= p3_tuple_8861_comb;
  end
  // __tmp__Butterfly_21___itok__tmp__Butterfly___itok__tmp__Butterfly_15___itok__apfloat__sub__8_23___itok__apfloat__sub__8_23_10___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p2_and_7971_comb | p2_and_7970_comb | p2_and_7969_comb)) p2_and_7971_comb | p2_and_7970_comb | p2_and_7969_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  // __tmp__Butterfly_21___itok__tmp__Butterfly___itok__tmp__Butterfly_16___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p2_and_7978_comb | p2_and_7977_comb | p2_and_7976_comb)) p2_and_7978_comb | p2_and_7977_comb | p2_and_7976_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  // __tmp__Butterfly_21___itok__tmp__Butterfly___itok__tmp__Butterfly_17___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p3_and_8497_comb | p3_and_8496_comb | p3_and_8495_comb)) p3_and_8497_comb | p3_and_8496_comb | p3_and_8495_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  // __tmp__Butterfly_21___itok__tmp__Butterfly___itok__tmp__Butterfly_18___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p3_and_8504_comb | p3_and_8503_comb | p3_and_8502_comb)) p3_and_8504_comb | p3_and_8503_comb | p3_and_8502_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  // __tmp__Butterfly_21___itok__tmp__Butterfly___itok__tmp__Butterfly_19___itok__apfloat__sub__8_23___itok__apfloat__sub__8_23_10___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p3_and_8511_comb | p3_and_8510_comb | p3_and_8509_comb)) p3_and_8511_comb | p3_and_8510_comb | p3_and_8509_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  // __tmp__Butterfly_21___itok__tmp__Butterfly___itok__tmp__Butterfly_20___itok__apfloat__sub__8_23___itok__apfloat__sub__8_23_10___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p3_and_8518_comb | p3_and_8517_comb | p3_and_8516_comb)) p3_and_8518_comb | p3_and_8517_comb | p3_and_8516_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  assign out = p3_tuple_8861;
endmodule
