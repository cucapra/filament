module Const #(
  parameter WIDTH = 32,
  parameter VALUE = 0
) (
  output wire logic [WIDTH-1:0] out
);
  assign out = VALUE;
endmodule

//// =========== Computation ============

module Add #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] left,
  input wire logic [IN_WIDTH-1:0] right,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module Sub #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] left,
  input wire logic [IN_WIDTH-1:0] right,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module MultComb #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] left,
  input wire logic [IN_WIDTH-1:0] right,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = left * right;
endmodule

//// =========== Binary Logical Operations ============

module And #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH-1:0] left,
  input wire logic [WIDTH-1:0] right,
  output wire logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module Or #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module Xor #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module Not #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] in,
  output wire logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

//// =========== Comparions ============

module Gt #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left > right;
endmodule

module Eq #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left == right;
endmodule

module Neq #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left != right;
endmodule

module Lt #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left < right;
endmodule

module Gte #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left >= right;
endmodule

module Lte #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left <= right;
endmodule

//// =========== Extension ============

module SignExtend #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  parameter EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = {{EXTEND{in[IN_WIDTH-1]}}, in};
endmodule

module ZeroExtend #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  parameter EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = {{EXTEND{1'b0}}, in};
endmodule

module Extend #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = {OUT_WIDTH{in}};
endmodule

module Concat #(
  parameter LEFT = 32,
  parameter RIGHT = 32,
  parameter OUT = 64
) (
  input wire logic [LEFT-1:0] left,
  input wire logic [RIGHT-1:0] right,
  output wire logic [OUT-1:0] out
);
  assign out = {left, right};
endmodule

//// =========== Select bits ============
module Select #(
  parameter WIDTH = 32,
  parameter POS = 0
) (
  input wire logic [WIDTH-1:0] in,
  output wire logic out
);
  assign out = in[POS];
endmodule

module Slice #(
  parameter IN_WIDTH = 32,
  parameter MSB = 31,
  parameter LSB = 0,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = in[MSB:LSB];
endmodule

/// =========== Reduction Operations ============
module ReduceAnd #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  output wire logic out
);
  assign out = &in;
endmodule

module ReduceOr #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  output wire logic out
);
  assign out = |in;
endmodule

/// ========== Shift Operations ============
module ShiftLeft #(
  parameter WIDTH = 32,
  parameter SHIFT_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  input wire logic [SHIFT_WIDTH-1:0] shift,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = in << shift;
endmodule

module ShiftRight #(
  parameter WIDTH = 32,
  parameter SHIFT_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  input wire logic [SHIFT_WIDTH-1:0] shift,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = in >> shift;
endmodule

module ArithShiftRight #(
  parameter WIDTH = 32
) (
  input wire logic signed [WIDTH-1:0] in,
  input wire logic [WIDTH-1:0] shift,
  output wire logic [WIDTH-1:0] out
); 
  assign out = in >>> shift;
endmodule

module Mux #(
  parameter WIDTH = 32
) (
  input wire logic sel,
  input wire logic [WIDTH-1:0] in0,
  input wire logic [WIDTH-1:0] in1,
  output logic [WIDTH-1:0] out
);
  assign out = sel ? in0 : in1;
endmodule
module Butterfly_Exp8_Mant23(
  input wire clk,
  input wire [31:0] in0_r,
  input wire [31:0] in0_i,
  input wire [31:0] in1_r,
  input wire [31:0] in1_i,
  input wire [31:0] twd_r,
  input wire [31:0] twd_i,
  output wire [127:0] out
);
  // lint_off MULTIPLY
  function automatic [47:0] umul48b_24b_x_24b (input reg [23:0] lhs, input reg [23:0] rhs);
    begin
      umul48b_24b_x_24b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_in0_r;
  reg [31:0] p0_in0_i;
  reg [31:0] p0_in1_r;
  reg [31:0] p0_in1_i;
  reg [31:0] p0_twd_r;
  reg [31:0] p0_twd_i;
  always_ff @ (posedge clk) begin
    p0_in0_r <= in0_r;
    p0_in0_i <= in0_i;
    p0_in1_r <= in1_r;
    p0_in1_i <= in1_i;
    p0_twd_r <= twd_r;
    p0_twd_i <= twd_i;
  end

  // ===== Pipe stage 1:
  wire [22:0] p1_in1_r_fraction__10_comb;
  wire [7:0] p1_in1_r_bexp__9_comb;
  wire [22:0] p1_twd_r_fraction__10_comb;
  wire [7:0] p1_twd_r_bexp__9_comb;
  wire [22:0] p1_in1_i_fraction__10_comb;
  wire [7:0] p1_in1_i_bexp__9_comb;
  wire [22:0] p1_twd_i_fraction__10_comb;
  wire [7:0] p1_twd_i_bexp__9_comb;
  wire [23:0] p1_in1_r_fraction__11_comb;
  wire [23:0] p1_twd_r_fraction__11_comb;
  wire [23:0] p1_in1_i_fraction__11_comb;
  wire [23:0] p1_twd_i_fraction__11_comb;
  wire [8:0] p1_concat_7295_comb;
  wire [8:0] p1_concat_7296_comb;
  wire [23:0] p1_in1_r_fraction__12_comb;
  wire [23:0] p1_twd_r_fraction__12_comb;
  wire [8:0] p1_concat_7301_comb;
  wire [8:0] p1_concat_7302_comb;
  wire [23:0] p1_in1_i_fraction__12_comb;
  wire [23:0] p1_twd_i_fraction__12_comb;
  wire [8:0] p1_add_7308_comb;
  wire p1_eq_7309_comb;
  wire p1_eq_7310_comb;
  wire [47:0] p1_fraction__1_comb;
  wire [8:0] p1_add_7313_comb;
  wire p1_eq_7314_comb;
  wire p1_eq_7315_comb;
  wire [47:0] p1_fraction__8_comb;
  wire [8:0] p1_add_7318_comb;
  wire [47:0] p1_fraction__16_comb;
  wire [8:0] p1_add_7321_comb;
  wire [47:0] p1_fraction__24_comb;
  wire [9:0] p1_exp__1_comb;
  wire [47:0] p1_fraction__2_comb;
  wire [47:0] p1_sticky__1_comb;
  wire [9:0] p1_exp__4_comb;
  wire [47:0] p1_fraction__9_comb;
  wire [47:0] p1_sticky__2_comb;
  wire [9:0] p1_exp__8_comb;
  wire [47:0] p1_fraction__17_comb;
  wire [47:0] p1_sticky__4_comb;
  wire [9:0] p1_exp__12_comb;
  wire [47:0] p1_fraction__25_comb;
  wire [47:0] p1_sticky__6_comb;
  wire [9:0] p1_exp__2_comb;
  wire [47:0] p1_fraction__3_comb;
  wire [9:0] p1_exp__5_comb;
  wire [47:0] p1_fraction__10_comb;
  wire [9:0] p1_exp__9_comb;
  wire [47:0] p1_fraction__18_comb;
  wire [9:0] p1_exp__13_comb;
  wire [47:0] p1_fraction__26_comb;
  wire [9:0] p1_exp__3_comb;
  wire [9:0] p1_exp__6_comb;
  wire [9:0] p1_exp__10_comb;
  wire [9:0] p1_exp__14_comb;
  wire [47:0] p1_fraction__4_comb;
  wire [47:0] p1_sticky__5_comb;
  wire [47:0] p1_fraction__11_comb;
  wire [47:0] p1_sticky__3_comb;
  wire [47:0] p1_fraction__19_comb;
  wire [47:0] p1_sticky__7_comb;
  wire [47:0] p1_fraction__27_comb;
  wire [47:0] p1_sticky__8_comb;
  wire [47:0] p1_fraction__5_comb;
  wire [47:0] p1_fraction__12_comb;
  wire [47:0] p1_fraction__20_comb;
  wire [47:0] p1_fraction__28_comb;
  wire [22:0] p1_fraction__6_comb;
  wire [22:0] p1_fraction__13_comb;
  wire [22:0] p1_fraction__21_comb;
  wire [22:0] p1_fraction__29_comb;
  wire p1_greater_than_half_way__2_comb;
  wire [23:0] p1_fraction__7_comb;
  wire p1_greater_than_half_way__1_comb;
  wire [23:0] p1_fraction__14_comb;
  wire p1_greater_than_half_way__3_comb;
  wire [23:0] p1_fraction__22_comb;
  wire p1_greater_than_half_way__4_comb;
  wire [23:0] p1_fraction__30_comb;
  wire p1_do_round_up__2_comb;
  wire [23:0] p1_add_7476_comb;
  wire p1_do_round_up__1_comb;
  wire [23:0] p1_add_7478_comb;
  wire p1_do_round_up__3_comb;
  wire [23:0] p1_add_7480_comb;
  wire p1_do_round_up__4_comb;
  wire [23:0] p1_add_7482_comb;
  wire [23:0] p1_fraction__23_comb;
  wire [23:0] p1_fraction__15_comb;
  wire [23:0] p1_fraction__31_comb;
  wire [23:0] p1_fraction__32_comb;
  wire [9:0] p1_add_7492_comb;
  wire [9:0] p1_add_7494_comb;
  wire [9:0] p1_add_7496_comb;
  wire [9:0] p1_add_7498_comb;
  wire [9:0] p1_exp__11_comb;
  wire [9:0] p1_exp__7_comb;
  wire [9:0] p1_exp__15_comb;
  wire [9:0] p1_exp__16_comb;
  wire p1_sgt_7507_comb;
  wire p1_sgt_7508_comb;
  wire p1_sgt_7509_comb;
  wire p1_sgt_7510_comb;
  wire [8:0] p1_result_exp__1_comb;
  wire [7:0] p1_high_exp__3_comb;
  wire [7:0] p1_high_exp__4_comb;
  wire [8:0] p1_result_exp__2_comb;
  wire [7:0] p1_high_exp__6_comb;
  wire [7:0] p1_high_exp__1_comb;
  wire [8:0] p1_result_exp__6_comb;
  wire [8:0] p1_result_exp__9_comb;
  wire [8:0] p1_result_exp__4_comb;
  wire p1_eq_7528_comb;
  wire p1_eq_7530_comb;
  wire [8:0] p1_result_exp__3_comb;
  wire p1_eq_7533_comb;
  wire p1_eq_7535_comb;
  wire [8:0] p1_result_exp__7_comb;
  wire [8:0] p1_result_exp__10_comb;
  wire p1_and_7549_comb;
  wire p1_and_7550_comb;
  wire p1_and_7561_comb;
  wire p1_and_7562_comb;
  wire p1_has_0_arg__2_comb;
  wire p1_has_inf_arg__2_comb;
  wire p1_has_0_arg__1_comb;
  wire p1_has_inf_arg__1_comb;
  wire p1_has_0_arg__3_comb;
  wire p1_has_inf_arg__3_comb;
  wire p1_has_0_arg__4_comb;
  wire p1_has_inf_arg__4_comb;
  wire p1_nor_7599_comb;
  wire p1_and_7601_comb;
  wire p1_and_7602_comb;
  wire p1_nor_7604_comb;
  wire p1_and_7606_comb;
  wire p1_and_7607_comb;
  wire p1_nor_7609_comb;
  wire p1_nor_7612_comb;
  wire [22:0] p1_result_fraction__3_comb;
  wire p1_is_result_nan__2_comb;
  wire [22:0] p1_result_fraction__1_comb;
  wire p1_is_result_nan__1_comb;
  wire [22:0] p1_result_fraction__6_comb;
  wire p1_is_result_nan__3_comb;
  wire [22:0] p1_result_fraction__9_comb;
  wire p1_is_result_nan__4_comb;
  wire [22:0] p1_result_fraction__4_comb;
  wire [22:0] p1_nan_fraction__1_comb;
  wire [7:0] p1_high_exp__29_comb;
  wire [22:0] p1_result_fraction__2_comb;
  wire [22:0] p1_nan_fraction__5_comb;
  wire [7:0] p1_high_exp__28_comb;
  wire [22:0] p1_result_fraction__7_comb;
  wire [22:0] p1_nan_fraction__3_comb;
  wire [7:0] p1_high_exp__30_comb;
  wire [22:0] p1_result_fraction__10_comb;
  wire [22:0] p1_nan_fraction__4_comb;
  wire [7:0] p1_high_exp__31_comb;
  wire [22:0] p1_result_fraction__8_comb;
  wire [7:0] p1_result_exp__8_comb;
  wire [22:0] p1_result_fraction__5_comb;
  wire [7:0] p1_result_exp__5_comb;
  wire [22:0] p1_result_fraction__11_comb;
  wire [7:0] p1_result_exp__11_comb;
  wire [22:0] p1_result_fraction__12_comb;
  wire [7:0] p1_result_exp__12_comb;
  wire [5:0] p1_add_7694_comb;
  wire p1_ugt_7696_comb;
  wire [5:0] p1_add_7700_comb;
  wire [5:0] p1_add_7705_comb;
  wire p1_ugt_7707_comb;
  wire [5:0] p1_add_7711_comb;
  wire [27:0] p1_wide_x_comb;
  wire [7:0] p1_greater_exp_bexp_comb;
  wire [27:0] p1_wide_y_comb;
  wire [27:0] p1_wide_x__2_comb;
  wire [7:0] p1_greater_exp_bexp__1_comb;
  wire [27:0] p1_wide_y__2_comb;
  wire [27:0] p1_wide_x__1_comb;
  wire [7:0] p1_sub_7728_comb;
  wire [27:0] p1_wide_y__1_comb;
  wire [7:0] p1_sub_7730_comb;
  wire [27:0] p1_wide_x__3_comb;
  wire [7:0] p1_sub_7732_comb;
  wire [27:0] p1_wide_y__3_comb;
  wire [7:0] p1_sub_7734_comb;
  wire p1_in1_i_sign__2_comb;
  wire p1_twd_i_sign__2_comb;
  wire [27:0] p1_dropped_x_comb;
  wire [27:0] p1_dropped_y_comb;
  wire [27:0] p1_dropped_x__1_comb;
  wire [27:0] p1_dropped_y__1_comb;
  wire p1_result_sign__2_comb;
  wire p1_in1_r_sign__2_comb;
  wire p1_twd_r_sign__2_comb;
  wire p1_result_sign__3_comb;
  wire p1_result_sign__1_comb;
  wire [7:0] p1_shift_x_comb;
  wire p1_sticky_x_comb;
  wire [7:0] p1_shift_y_comb;
  wire p1_sticky_y_comb;
  wire p1_result_sign__6_comb;
  wire p1_result_sign__4_comb;
  wire [7:0] p1_shift_x__1_comb;
  wire p1_sticky_x__1_comb;
  wire [7:0] p1_shift_y__1_comb;
  wire p1_sticky_y__1_comb;
  wire p1_bd__1_sign_comb;
  wire p1_result_sign__5_comb;
  wire [27:0] p1_shifted_x_comb;
  wire [27:0] p1_shifted_y_comb;
  wire p1_result_sign__8_comb;
  wire p1_result_sign__7_comb;
  wire [27:0] p1_shifted_x__1_comb;
  wire [27:0] p1_shifted_y__1_comb;
  wire [7:0] p1_high_exp__32_comb;
  wire [7:0] p1_high_exp__33_comb;
  wire [7:0] p1_high_exp__34_comb;
  wire [7:0] p1_high_exp__35_comb;
  wire p1_greater_exp_sign_comb;
  wire [27:0] p1_addend_x_comb;
  wire [27:0] p1_addend_y_comb;
  wire p1_greater_exp_sign__1_comb;
  wire [27:0] p1_addend_x__2_comb;
  wire [27:0] p1_addend_y__2_comb;
  wire p1_eq_7824_comb;
  wire p1_eq_7825_comb;
  wire p1_eq_7826_comb;
  wire p1_eq_7827_comb;
  wire p1_eq_7828_comb;
  wire p1_eq_7829_comb;
  wire p1_eq_7830_comb;
  wire p1_eq_7831_comb;
  wire p1_and_7834_comb;
  wire p1_and_7835_comb;
  wire p1_and_7838_comb;
  wire p1_and_7839_comb;
  wire [27:0] p1_addend_x__1_comb;
  wire [27:0] p1_addend_y__1_comb;
  wire [27:0] p1_addend_x__3_comb;
  wire [27:0] p1_addend_y__3_comb;
  wire p1_has_pos_inf_comb;
  wire p1_has_neg_inf_comb;
  wire p1_has_pos_inf__1_comb;
  wire p1_has_neg_inf__1_comb;
  wire [28:0] p1_fraction__33_comb;
  wire [28:0] p1_fraction__34_comb;
  wire [27:0] p1_bit_slice_7808_comb;
  wire [27:0] p1_bit_slice_7809_comb;
  wire p1_bit_slice_7810_comb;
  wire p1_bit_slice_7811_comb;
  wire p1_ne_7814_comb;
  wire p1_ne_7815_comb;
  wire p1_nor_7860_comb;
  wire p1_nor_7864_comb;
  wire p1_is_result_nan__5_comb;
  wire p1_is_operand_inf_comb;
  wire p1_is_result_nan__6_comb;
  wire p1_is_operand_inf__1_comb;
  wire [22:0] p1_in0_r_fraction__6_comb;
  wire [7:0] p1_in0_r_bexp__6_comb;
  wire [22:0] p1_in0_i_fraction__6_comb;
  wire [7:0] p1_in0_i_bexp__6_comb;
  wire p1_fraction_is_zero_comb;
  wire p1_fraction_is_zero__1_comb;
  wire p1_not_7880_comb;
  wire p1_not_7881_comb;
  wire p1_in0_r_sign__2_comb;
  wire p1_in0_i_sign__2_comb;
  assign p1_in1_r_fraction__10_comb = p0_in1_r[22:0];
  assign p1_in1_r_bexp__9_comb = p0_in1_r[30:23];
  assign p1_twd_r_fraction__10_comb = p0_twd_r[22:0];
  assign p1_twd_r_bexp__9_comb = p0_twd_r[30:23];
  assign p1_in1_i_fraction__10_comb = p0_in1_i[22:0];
  assign p1_in1_i_bexp__9_comb = p0_in1_i[30:23];
  assign p1_twd_i_fraction__10_comb = p0_twd_i[22:0];
  assign p1_twd_i_bexp__9_comb = p0_twd_i[30:23];
  assign p1_in1_r_fraction__11_comb = {1'h0, p1_in1_r_fraction__10_comb} | 24'h80_0000;
  assign p1_twd_r_fraction__11_comb = {1'h0, p1_twd_r_fraction__10_comb} | 24'h80_0000;
  assign p1_in1_i_fraction__11_comb = {1'h0, p1_in1_i_fraction__10_comb} | 24'h80_0000;
  assign p1_twd_i_fraction__11_comb = {1'h0, p1_twd_i_fraction__10_comb} | 24'h80_0000;
  assign p1_concat_7295_comb = {1'h0, p1_in1_r_bexp__9_comb};
  assign p1_concat_7296_comb = {1'h0, p1_twd_r_bexp__9_comb};
  assign p1_in1_r_fraction__12_comb = p1_in1_r_fraction__11_comb & {24{p1_in1_r_bexp__9_comb != 8'h00}};
  assign p1_twd_r_fraction__12_comb = p1_twd_r_fraction__11_comb & {24{p1_twd_r_bexp__9_comb != 8'h00}};
  assign p1_concat_7301_comb = {1'h0, p1_in1_i_bexp__9_comb};
  assign p1_concat_7302_comb = {1'h0, p1_twd_i_bexp__9_comb};
  assign p1_in1_i_fraction__12_comb = p1_in1_i_fraction__11_comb & {24{p1_in1_i_bexp__9_comb != 8'h00}};
  assign p1_twd_i_fraction__12_comb = p1_twd_i_fraction__11_comb & {24{p1_twd_i_bexp__9_comb != 8'h00}};
  assign p1_add_7308_comb = p1_concat_7295_comb + p1_concat_7296_comb;
  assign p1_eq_7309_comb = p1_in1_r_bexp__9_comb == 8'h00;
  assign p1_eq_7310_comb = p1_twd_r_bexp__9_comb == 8'h00;
  assign p1_fraction__1_comb = umul48b_24b_x_24b(p1_in1_r_fraction__12_comb, p1_twd_r_fraction__12_comb);
  assign p1_add_7313_comb = p1_concat_7301_comb + p1_concat_7302_comb;
  assign p1_eq_7314_comb = p1_in1_i_bexp__9_comb == 8'h00;
  assign p1_eq_7315_comb = p1_twd_i_bexp__9_comb == 8'h00;
  assign p1_fraction__8_comb = umul48b_24b_x_24b(p1_in1_i_fraction__12_comb, p1_twd_i_fraction__12_comb);
  assign p1_add_7318_comb = p1_concat_7295_comb + p1_concat_7302_comb;
  assign p1_fraction__16_comb = umul48b_24b_x_24b(p1_in1_r_fraction__12_comb, p1_twd_i_fraction__12_comb);
  assign p1_add_7321_comb = p1_concat_7301_comb + p1_concat_7296_comb;
  assign p1_fraction__24_comb = umul48b_24b_x_24b(p1_in1_i_fraction__12_comb, p1_twd_r_fraction__12_comb);
  assign p1_exp__1_comb = {1'h0, p1_add_7308_comb} + 10'h381;
  assign p1_fraction__2_comb = p1_fraction__1_comb >> p1_fraction__1_comb[47];
  assign p1_sticky__1_comb = {47'h0000_0000_0000, p1_fraction__1_comb[0]};
  assign p1_exp__4_comb = {1'h0, p1_add_7313_comb} + 10'h381;
  assign p1_fraction__9_comb = p1_fraction__8_comb >> p1_fraction__8_comb[47];
  assign p1_sticky__2_comb = {47'h0000_0000_0000, p1_fraction__8_comb[0]};
  assign p1_exp__8_comb = {1'h0, p1_add_7318_comb} + 10'h381;
  assign p1_fraction__17_comb = p1_fraction__16_comb >> p1_fraction__16_comb[47];
  assign p1_sticky__4_comb = {47'h0000_0000_0000, p1_fraction__16_comb[0]};
  assign p1_exp__12_comb = {1'h0, p1_add_7321_comb} + 10'h381;
  assign p1_fraction__25_comb = p1_fraction__24_comb >> p1_fraction__24_comb[47];
  assign p1_sticky__6_comb = {47'h0000_0000_0000, p1_fraction__24_comb[0]};
  assign p1_exp__2_comb = p1_exp__1_comb & {10{~(p1_eq_7309_comb | p1_eq_7310_comb)}};
  assign p1_fraction__3_comb = p1_fraction__2_comb | p1_sticky__1_comb;
  assign p1_exp__5_comb = p1_exp__4_comb & {10{~(p1_eq_7314_comb | p1_eq_7315_comb)}};
  assign p1_fraction__10_comb = p1_fraction__9_comb | p1_sticky__2_comb;
  assign p1_exp__9_comb = p1_exp__8_comb & {10{~(p1_eq_7309_comb | p1_eq_7315_comb)}};
  assign p1_fraction__18_comb = p1_fraction__17_comb | p1_sticky__4_comb;
  assign p1_exp__13_comb = p1_exp__12_comb & {10{~(p1_eq_7314_comb | p1_eq_7310_comb)}};
  assign p1_fraction__26_comb = p1_fraction__25_comb | p1_sticky__6_comb;
  assign p1_exp__3_comb = p1_exp__2_comb + {9'h000, p1_fraction__1_comb[47]};
  assign p1_exp__6_comb = p1_exp__5_comb + {9'h000, p1_fraction__8_comb[47]};
  assign p1_exp__10_comb = p1_exp__9_comb + {9'h000, p1_fraction__16_comb[47]};
  assign p1_exp__14_comb = p1_exp__13_comb + {9'h000, p1_fraction__24_comb[47]};
  assign p1_fraction__4_comb = $signed(p1_exp__3_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__3_comb[47:1]} : p1_fraction__3_comb;
  assign p1_sticky__5_comb = {47'h0000_0000_0000, p1_fraction__3_comb[0]};
  assign p1_fraction__11_comb = $signed(p1_exp__6_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__10_comb[47:1]} : p1_fraction__10_comb;
  assign p1_sticky__3_comb = {47'h0000_0000_0000, p1_fraction__10_comb[0]};
  assign p1_fraction__19_comb = $signed(p1_exp__10_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__18_comb[47:1]} : p1_fraction__18_comb;
  assign p1_sticky__7_comb = {47'h0000_0000_0000, p1_fraction__18_comb[0]};
  assign p1_fraction__27_comb = $signed(p1_exp__14_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__26_comb[47:1]} : p1_fraction__26_comb;
  assign p1_sticky__8_comb = {47'h0000_0000_0000, p1_fraction__26_comb[0]};
  assign p1_fraction__5_comb = p1_fraction__4_comb | p1_sticky__5_comb;
  assign p1_fraction__12_comb = p1_fraction__11_comb | p1_sticky__3_comb;
  assign p1_fraction__20_comb = p1_fraction__19_comb | p1_sticky__7_comb;
  assign p1_fraction__28_comb = p1_fraction__27_comb | p1_sticky__8_comb;
  assign p1_fraction__6_comb = p1_fraction__5_comb[45:23];
  assign p1_fraction__13_comb = p1_fraction__12_comb[45:23];
  assign p1_fraction__21_comb = p1_fraction__20_comb[45:23];
  assign p1_fraction__29_comb = p1_fraction__28_comb[45:23];
  assign p1_greater_than_half_way__2_comb = p1_fraction__5_comb[22] & p1_fraction__5_comb[21:0] != 22'h00_0000;
  assign p1_fraction__7_comb = {1'h0, p1_fraction__6_comb};
  assign p1_greater_than_half_way__1_comb = p1_fraction__12_comb[22] & p1_fraction__12_comb[21:0] != 22'h00_0000;
  assign p1_fraction__14_comb = {1'h0, p1_fraction__13_comb};
  assign p1_greater_than_half_way__3_comb = p1_fraction__20_comb[22] & p1_fraction__20_comb[21:0] != 22'h00_0000;
  assign p1_fraction__22_comb = {1'h0, p1_fraction__21_comb};
  assign p1_greater_than_half_way__4_comb = p1_fraction__28_comb[22] & p1_fraction__28_comb[21:0] != 22'h00_0000;
  assign p1_fraction__30_comb = {1'h0, p1_fraction__29_comb};
  assign p1_do_round_up__2_comb = p1_greater_than_half_way__2_comb | p1_fraction__5_comb[22] & p1_fraction__5_comb[21:0] == 22'h00_0000 & p1_fraction__5_comb[23];
  assign p1_add_7476_comb = p1_fraction__7_comb + 24'h00_0001;
  assign p1_do_round_up__1_comb = p1_greater_than_half_way__1_comb | p1_fraction__12_comb[22] & p1_fraction__12_comb[21:0] == 22'h00_0000 & p1_fraction__12_comb[23];
  assign p1_add_7478_comb = p1_fraction__14_comb + 24'h00_0001;
  assign p1_do_round_up__3_comb = p1_greater_than_half_way__3_comb | p1_fraction__20_comb[22] & p1_fraction__20_comb[21:0] == 22'h00_0000 & p1_fraction__20_comb[23];
  assign p1_add_7480_comb = p1_fraction__22_comb + 24'h00_0001;
  assign p1_do_round_up__4_comb = p1_greater_than_half_way__4_comb | p1_fraction__28_comb[22] & p1_fraction__28_comb[21:0] == 22'h00_0000 & p1_fraction__28_comb[23];
  assign p1_add_7482_comb = p1_fraction__30_comb + 24'h00_0001;
  assign p1_fraction__23_comb = p1_do_round_up__2_comb ? p1_add_7476_comb : p1_fraction__7_comb;
  assign p1_fraction__15_comb = p1_do_round_up__1_comb ? p1_add_7478_comb : p1_fraction__14_comb;
  assign p1_fraction__31_comb = p1_do_round_up__3_comb ? p1_add_7480_comb : p1_fraction__22_comb;
  assign p1_fraction__32_comb = p1_do_round_up__4_comb ? p1_add_7482_comb : p1_fraction__30_comb;
  assign p1_add_7492_comb = p1_exp__3_comb + 10'h001;
  assign p1_add_7494_comb = p1_exp__6_comb + 10'h001;
  assign p1_add_7496_comb = p1_exp__10_comb + 10'h001;
  assign p1_add_7498_comb = p1_exp__14_comb + 10'h001;
  assign p1_exp__11_comb = p1_fraction__23_comb[23] ? p1_add_7492_comb : p1_exp__3_comb;
  assign p1_exp__7_comb = p1_fraction__15_comb[23] ? p1_add_7494_comb : p1_exp__6_comb;
  assign p1_exp__15_comb = p1_fraction__31_comb[23] ? p1_add_7496_comb : p1_exp__10_comb;
  assign p1_exp__16_comb = p1_fraction__32_comb[23] ? p1_add_7498_comb : p1_exp__14_comb;
  assign p1_sgt_7507_comb = $signed(p1_exp__11_comb) > $signed(10'h000);
  assign p1_sgt_7508_comb = $signed(p1_exp__7_comb) > $signed(10'h000);
  assign p1_sgt_7509_comb = $signed(p1_exp__15_comb) > $signed(10'h000);
  assign p1_sgt_7510_comb = $signed(p1_exp__16_comb) > $signed(10'h000);
  assign p1_result_exp__1_comb = p1_exp__11_comb[8:0];
  assign p1_high_exp__3_comb = 8'hff;
  assign p1_high_exp__4_comb = 8'hff;
  assign p1_result_exp__2_comb = p1_exp__7_comb[8:0];
  assign p1_high_exp__6_comb = 8'hff;
  assign p1_high_exp__1_comb = 8'hff;
  assign p1_result_exp__6_comb = p1_exp__15_comb[8:0];
  assign p1_result_exp__9_comb = p1_exp__16_comb[8:0];
  assign p1_result_exp__4_comb = p1_result_exp__1_comb & {9{p1_sgt_7507_comb}};
  assign p1_eq_7528_comb = p1_in1_r_bexp__9_comb == p1_high_exp__3_comb;
  assign p1_eq_7530_comb = p1_twd_r_bexp__9_comb == p1_high_exp__4_comb;
  assign p1_result_exp__3_comb = p1_result_exp__2_comb & {9{p1_sgt_7508_comb}};
  assign p1_eq_7533_comb = p1_in1_i_bexp__9_comb == p1_high_exp__6_comb;
  assign p1_eq_7535_comb = p1_twd_i_bexp__9_comb == p1_high_exp__1_comb;
  assign p1_result_exp__7_comb = p1_result_exp__6_comb & {9{p1_sgt_7509_comb}};
  assign p1_result_exp__10_comb = p1_result_exp__9_comb & {9{p1_sgt_7510_comb}};
  assign p1_and_7549_comb = p1_eq_7528_comb & p1_in1_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_7550_comb = p1_eq_7530_comb & p1_twd_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_7561_comb = p1_eq_7533_comb & p1_in1_i_fraction__10_comb == 23'h00_0000;
  assign p1_and_7562_comb = p1_eq_7535_comb & p1_twd_i_fraction__10_comb == 23'h00_0000;
  assign p1_has_0_arg__2_comb = p1_eq_7309_comb | p1_eq_7310_comb;
  assign p1_has_inf_arg__2_comb = p1_and_7549_comb | p1_and_7550_comb;
  assign p1_has_0_arg__1_comb = p1_eq_7314_comb | p1_eq_7315_comb;
  assign p1_has_inf_arg__1_comb = p1_and_7561_comb | p1_and_7562_comb;
  assign p1_has_0_arg__3_comb = p1_eq_7309_comb | p1_eq_7315_comb;
  assign p1_has_inf_arg__3_comb = p1_and_7549_comb | p1_and_7562_comb;
  assign p1_has_0_arg__4_comb = p1_eq_7314_comb | p1_eq_7310_comb;
  assign p1_has_inf_arg__4_comb = p1_and_7561_comb | p1_and_7550_comb;
  assign p1_nor_7599_comb = ~(p1_result_exp__4_comb[8] | p1_result_exp__4_comb[0] & p1_result_exp__4_comb[1] & p1_result_exp__4_comb[2] & p1_result_exp__4_comb[3] & p1_result_exp__4_comb[4] & p1_result_exp__4_comb[5] & p1_result_exp__4_comb[6] & p1_result_exp__4_comb[7]);
  assign p1_and_7601_comb = p1_eq_7528_comb & p1_in1_r_fraction__10_comb != 23'h00_0000;
  assign p1_and_7602_comb = p1_eq_7530_comb & p1_twd_r_fraction__10_comb != 23'h00_0000;
  assign p1_nor_7604_comb = ~(p1_result_exp__3_comb[8] | p1_result_exp__3_comb[0] & p1_result_exp__3_comb[1] & p1_result_exp__3_comb[2] & p1_result_exp__3_comb[3] & p1_result_exp__3_comb[4] & p1_result_exp__3_comb[5] & p1_result_exp__3_comb[6] & p1_result_exp__3_comb[7]);
  assign p1_and_7606_comb = p1_eq_7533_comb & p1_in1_i_fraction__10_comb != 23'h00_0000;
  assign p1_and_7607_comb = p1_eq_7535_comb & p1_twd_i_fraction__10_comb != 23'h00_0000;
  assign p1_nor_7609_comb = ~(p1_result_exp__7_comb[8] | p1_result_exp__7_comb[0] & p1_result_exp__7_comb[1] & p1_result_exp__7_comb[2] & p1_result_exp__7_comb[3] & p1_result_exp__7_comb[4] & p1_result_exp__7_comb[5] & p1_result_exp__7_comb[6] & p1_result_exp__7_comb[7]);
  assign p1_nor_7612_comb = ~(p1_result_exp__10_comb[8] | p1_result_exp__10_comb[0] & p1_result_exp__10_comb[1] & p1_result_exp__10_comb[2] & p1_result_exp__10_comb[3] & p1_result_exp__10_comb[4] & p1_result_exp__10_comb[5] & p1_result_exp__10_comb[6] & p1_result_exp__10_comb[7]);
  assign p1_result_fraction__3_comb = p1_fraction__23_comb[22:0];
  assign p1_is_result_nan__2_comb = p1_and_7601_comb | p1_and_7602_comb | p1_has_0_arg__2_comb & p1_has_inf_arg__2_comb;
  assign p1_result_fraction__1_comb = p1_fraction__15_comb[22:0];
  assign p1_is_result_nan__1_comb = p1_and_7606_comb | p1_and_7607_comb | p1_has_0_arg__1_comb & p1_has_inf_arg__1_comb;
  assign p1_result_fraction__6_comb = p1_fraction__31_comb[22:0];
  assign p1_is_result_nan__3_comb = p1_and_7601_comb | p1_and_7607_comb | p1_has_0_arg__3_comb & p1_has_inf_arg__3_comb;
  assign p1_result_fraction__9_comb = p1_fraction__32_comb[22:0];
  assign p1_is_result_nan__4_comb = p1_and_7606_comb | p1_and_7602_comb | p1_has_0_arg__4_comb & p1_has_inf_arg__4_comb;
  assign p1_result_fraction__4_comb = p1_result_fraction__3_comb & {23{p1_sgt_7507_comb}} & {23{p1_nor_7599_comb}} & {23{~(p1_and_7549_comb | p1_and_7550_comb)}};
  assign p1_nan_fraction__1_comb = 23'h40_0000;
  assign p1_high_exp__29_comb = 8'hff;
  assign p1_result_fraction__2_comb = p1_result_fraction__1_comb & {23{p1_sgt_7508_comb}} & {23{p1_nor_7604_comb}} & {23{~(p1_and_7561_comb | p1_and_7562_comb)}};
  assign p1_nan_fraction__5_comb = 23'h40_0000;
  assign p1_high_exp__28_comb = 8'hff;
  assign p1_result_fraction__7_comb = p1_result_fraction__6_comb & {23{p1_sgt_7509_comb}} & {23{p1_nor_7609_comb}} & {23{~(p1_and_7549_comb | p1_and_7562_comb)}};
  assign p1_nan_fraction__3_comb = 23'h40_0000;
  assign p1_high_exp__30_comb = 8'hff;
  assign p1_result_fraction__10_comb = p1_result_fraction__9_comb & {23{p1_sgt_7510_comb}} & {23{p1_nor_7612_comb}} & {23{~(p1_and_7561_comb | p1_and_7550_comb)}};
  assign p1_nan_fraction__4_comb = 23'h40_0000;
  assign p1_high_exp__31_comb = 8'hff;
  assign p1_result_fraction__8_comb = p1_is_result_nan__2_comb ? p1_nan_fraction__1_comb : p1_result_fraction__4_comb;
  assign p1_result_exp__8_comb = p1_is_result_nan__2_comb | p1_has_inf_arg__2_comb | ~p1_nor_7599_comb ? p1_high_exp__29_comb : p1_result_exp__4_comb[7:0];
  assign p1_result_fraction__5_comb = p1_is_result_nan__1_comb ? p1_nan_fraction__5_comb : p1_result_fraction__2_comb;
  assign p1_result_exp__5_comb = p1_is_result_nan__1_comb | p1_has_inf_arg__1_comb | ~p1_nor_7604_comb ? p1_high_exp__28_comb : p1_result_exp__3_comb[7:0];
  assign p1_result_fraction__11_comb = p1_is_result_nan__3_comb ? p1_nan_fraction__3_comb : p1_result_fraction__7_comb;
  assign p1_result_exp__11_comb = p1_is_result_nan__3_comb | p1_has_inf_arg__3_comb | ~p1_nor_7609_comb ? p1_high_exp__30_comb : p1_result_exp__7_comb[7:0];
  assign p1_result_fraction__12_comb = p1_is_result_nan__4_comb ? p1_nan_fraction__4_comb : p1_result_fraction__10_comb;
  assign p1_result_exp__12_comb = p1_is_result_nan__4_comb | p1_has_inf_arg__4_comb | ~p1_nor_7612_comb ? p1_high_exp__31_comb : p1_result_exp__10_comb[7:0];
  assign p1_add_7694_comb = p1_result_exp__8_comb[7:2] + 6'h07;
  assign p1_ugt_7696_comb = p1_result_exp__8_comb > p1_result_exp__5_comb;
  assign p1_add_7700_comb = p1_result_exp__5_comb[7:2] + 6'h07;
  assign p1_add_7705_comb = p1_result_exp__11_comb[7:2] + 6'h07;
  assign p1_ugt_7707_comb = p1_result_exp__11_comb > p1_result_exp__12_comb;
  assign p1_add_7711_comb = p1_result_exp__12_comb[7:2] + 6'h07;
  assign p1_wide_x_comb = {{2'h0, p1_result_fraction__8_comb} | 25'h080_0000, 3'h0};
  assign p1_greater_exp_bexp_comb = p1_ugt_7696_comb ? p1_result_exp__8_comb : p1_result_exp__5_comb;
  assign p1_wide_y_comb = {{2'h0, p1_result_fraction__5_comb} | 25'h080_0000, 3'h0};
  assign p1_wide_x__2_comb = {{2'h0, p1_result_fraction__11_comb} | 25'h080_0000, 3'h0};
  assign p1_greater_exp_bexp__1_comb = p1_ugt_7707_comb ? p1_result_exp__11_comb : p1_result_exp__12_comb;
  assign p1_wide_y__2_comb = {{2'h0, p1_result_fraction__12_comb} | 25'h080_0000, 3'h0};
  assign p1_wide_x__1_comb = p1_wide_x_comb & {28{p1_result_exp__8_comb != 8'h00}};
  assign p1_sub_7728_comb = {p1_add_7694_comb, p1_result_exp__8_comb[1:0]} - p1_greater_exp_bexp_comb;
  assign p1_wide_y__1_comb = p1_wide_y_comb & {28{p1_result_exp__5_comb != 8'h00}};
  assign p1_sub_7730_comb = {p1_add_7700_comb, p1_result_exp__5_comb[1:0]} - p1_greater_exp_bexp_comb;
  assign p1_wide_x__3_comb = p1_wide_x__2_comb & {28{p1_result_exp__11_comb != 8'h00}};
  assign p1_sub_7732_comb = {p1_add_7705_comb, p1_result_exp__11_comb[1:0]} - p1_greater_exp_bexp__1_comb;
  assign p1_wide_y__3_comb = p1_wide_y__2_comb & {28{p1_result_exp__12_comb != 8'h00}};
  assign p1_sub_7734_comb = {p1_add_7711_comb, p1_result_exp__12_comb[1:0]} - p1_greater_exp_bexp__1_comb;
  assign p1_in1_i_sign__2_comb = p0_in1_i[31:31];
  assign p1_twd_i_sign__2_comb = p0_twd_i[31:31];
  assign p1_dropped_x_comb = p1_sub_7728_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__1_comb << p1_sub_7728_comb;
  assign p1_dropped_y_comb = p1_sub_7730_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__1_comb << p1_sub_7730_comb;
  assign p1_dropped_x__1_comb = p1_sub_7732_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__3_comb << p1_sub_7732_comb;
  assign p1_dropped_y__1_comb = p1_sub_7734_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__3_comb << p1_sub_7734_comb;
  assign p1_result_sign__2_comb = p1_in1_i_sign__2_comb ^ p1_twd_i_sign__2_comb;
  assign p1_in1_r_sign__2_comb = p0_in1_r[31:31];
  assign p1_twd_r_sign__2_comb = p0_twd_r[31:31];
  assign p1_result_sign__3_comb = ~p1_is_result_nan__1_comb & p1_result_sign__2_comb;
  assign p1_result_sign__1_comb = p1_in1_r_sign__2_comb ^ p1_twd_r_sign__2_comb;
  assign p1_shift_x_comb = p1_greater_exp_bexp_comb - p1_result_exp__8_comb;
  assign p1_sticky_x_comb = p1_dropped_x_comb[27:3] != 25'h000_0000;
  assign p1_shift_y_comb = p1_greater_exp_bexp_comb - p1_result_exp__5_comb;
  assign p1_sticky_y_comb = p1_dropped_y_comb[27:3] != 25'h000_0000;
  assign p1_result_sign__6_comb = p1_in1_i_sign__2_comb ^ p1_twd_r_sign__2_comb;
  assign p1_result_sign__4_comb = p1_in1_r_sign__2_comb ^ p1_twd_i_sign__2_comb;
  assign p1_shift_x__1_comb = p1_greater_exp_bexp__1_comb - p1_result_exp__11_comb;
  assign p1_sticky_x__1_comb = p1_dropped_x__1_comb[27:3] != 25'h000_0000;
  assign p1_shift_y__1_comb = p1_greater_exp_bexp__1_comb - p1_result_exp__12_comb;
  assign p1_sticky_y__1_comb = p1_dropped_y__1_comb[27:3] != 25'h000_0000;
  assign p1_bd__1_sign_comb = ~p1_result_sign__3_comb;
  assign p1_result_sign__5_comb = ~p1_is_result_nan__2_comb & p1_result_sign__1_comb;
  assign p1_shifted_x_comb = p1_shift_x_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__1_comb >> p1_shift_x_comb;
  assign p1_shifted_y_comb = p1_shift_y_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__1_comb >> p1_shift_y_comb;
  assign p1_result_sign__8_comb = ~p1_is_result_nan__4_comb & p1_result_sign__6_comb;
  assign p1_result_sign__7_comb = ~p1_is_result_nan__3_comb & p1_result_sign__4_comb;
  assign p1_shifted_x__1_comb = p1_shift_x__1_comb >= 8'h1c ? 28'h000_0000 : p1_wide_x__3_comb >> p1_shift_x__1_comb;
  assign p1_shifted_y__1_comb = p1_shift_y__1_comb >= 8'h1c ? 28'h000_0000 : p1_wide_y__3_comb >> p1_shift_y__1_comb;
  assign p1_high_exp__32_comb = 8'hff;
  assign p1_high_exp__33_comb = 8'hff;
  assign p1_high_exp__34_comb = 8'hff;
  assign p1_high_exp__35_comb = 8'hff;
  assign p1_greater_exp_sign_comb = p1_ugt_7696_comb ? p1_result_sign__5_comb : p1_bd__1_sign_comb;
  assign p1_addend_x_comb = p1_shifted_x_comb | {27'h000_0000, p1_sticky_x_comb};
  assign p1_addend_y_comb = p1_shifted_y_comb | {27'h000_0000, p1_sticky_y_comb};
  assign p1_greater_exp_sign__1_comb = p1_ugt_7707_comb ? p1_result_sign__7_comb : p1_result_sign__8_comb;
  assign p1_addend_x__2_comb = p1_shifted_x__1_comb | {27'h000_0000, p1_sticky_x__1_comb};
  assign p1_addend_y__2_comb = p1_shifted_y__1_comb | {27'h000_0000, p1_sticky_y__1_comb};
  assign p1_eq_7824_comb = p1_result_exp__8_comb == p1_high_exp__32_comb;
  assign p1_eq_7825_comb = p1_result_fraction__8_comb == 23'h00_0000;
  assign p1_eq_7826_comb = p1_result_exp__5_comb == p1_high_exp__33_comb;
  assign p1_eq_7827_comb = p1_result_fraction__5_comb == 23'h00_0000;
  assign p1_eq_7828_comb = p1_result_exp__11_comb == p1_high_exp__34_comb;
  assign p1_eq_7829_comb = p1_result_fraction__11_comb == 23'h00_0000;
  assign p1_eq_7830_comb = p1_result_exp__12_comb == p1_high_exp__35_comb;
  assign p1_eq_7831_comb = p1_result_fraction__12_comb == 23'h00_0000;
  assign p1_and_7834_comb = p1_eq_7824_comb & p1_eq_7825_comb;
  assign p1_and_7835_comb = p1_eq_7826_comb & p1_eq_7827_comb;
  assign p1_and_7838_comb = p1_eq_7828_comb & p1_eq_7829_comb;
  assign p1_and_7839_comb = p1_eq_7830_comb & p1_eq_7831_comb;
  assign p1_addend_x__1_comb = p1_result_sign__5_comb ^ p1_greater_exp_sign_comb ? -p1_addend_x_comb : p1_addend_x_comb;
  assign p1_addend_y__1_comb = p1_bd__1_sign_comb ^ p1_greater_exp_sign_comb ? -p1_addend_y_comb : p1_addend_y_comb;
  assign p1_addend_x__3_comb = p1_result_sign__7_comb ^ p1_greater_exp_sign__1_comb ? -p1_addend_x__2_comb : p1_addend_x__2_comb;
  assign p1_addend_y__3_comb = p1_result_sign__8_comb ^ p1_greater_exp_sign__1_comb ? -p1_addend_y__2_comb : p1_addend_y__2_comb;
  assign p1_has_pos_inf_comb = ~(~(p1_eq_7824_comb & p1_eq_7825_comb) | p1_result_sign__5_comb) | ~(~(p1_eq_7826_comb & p1_eq_7827_comb) | p1_bd__1_sign_comb);
  assign p1_has_neg_inf_comb = p1_and_7834_comb & p1_result_sign__5_comb | p1_and_7835_comb & p1_bd__1_sign_comb;
  assign p1_has_pos_inf__1_comb = ~(~(p1_eq_7828_comb & p1_eq_7829_comb) | p1_result_sign__7_comb) | ~(~(p1_eq_7830_comb & p1_eq_7831_comb) | p1_result_sign__8_comb);
  assign p1_has_neg_inf__1_comb = p1_and_7838_comb & p1_result_sign__7_comb | p1_and_7839_comb & p1_result_sign__8_comb;
  assign p1_fraction__33_comb = {{1{p1_addend_x__1_comb[27]}}, p1_addend_x__1_comb} + {{1{p1_addend_y__1_comb[27]}}, p1_addend_y__1_comb};
  assign p1_fraction__34_comb = {{1{p1_addend_x__3_comb[27]}}, p1_addend_x__3_comb} + {{1{p1_addend_y__3_comb[27]}}, p1_addend_y__3_comb};
  assign p1_bit_slice_7808_comb = p1_fraction__33_comb[27:0];
  assign p1_bit_slice_7809_comb = p1_fraction__34_comb[27:0];
  assign p1_bit_slice_7810_comb = p1_fraction__33_comb[28];
  assign p1_bit_slice_7811_comb = p1_fraction__34_comb[28];
  assign p1_ne_7814_comb = p1_fraction__33_comb != 29'h0000_0000;
  assign p1_ne_7815_comb = p1_fraction__34_comb != 29'h0000_0000;
  assign p1_nor_7860_comb = ~(p1_and_7834_comb | p1_and_7835_comb);
  assign p1_nor_7864_comb = ~(p1_and_7838_comb | p1_and_7839_comb);
  assign p1_is_result_nan__5_comb = p1_eq_7824_comb & p1_result_fraction__8_comb != 23'h00_0000 | p1_eq_7826_comb & p1_result_fraction__5_comb != 23'h00_0000 | p1_has_pos_inf_comb & p1_has_neg_inf_comb;
  assign p1_is_operand_inf_comb = p1_and_7834_comb | p1_and_7835_comb;
  assign p1_is_result_nan__6_comb = p1_eq_7828_comb & p1_result_fraction__11_comb != 23'h00_0000 | p1_eq_7830_comb & p1_result_fraction__12_comb != 23'h00_0000 | p1_has_pos_inf__1_comb & p1_has_neg_inf__1_comb;
  assign p1_is_operand_inf__1_comb = p1_and_7838_comb | p1_and_7839_comb;
  assign p1_in0_r_fraction__6_comb = p0_in0_r[22:0];
  assign p1_in0_r_bexp__6_comb = p0_in0_r[30:23];
  assign p1_in0_i_fraction__6_comb = p0_in0_i[22:0];
  assign p1_in0_i_bexp__6_comb = p0_in0_i[30:23];
  assign p1_fraction_is_zero_comb = p1_fraction__33_comb == 29'h0000_0000;
  assign p1_fraction_is_zero__1_comb = p1_fraction__34_comb == 29'h0000_0000;
  assign p1_not_7880_comb = ~p1_has_pos_inf_comb;
  assign p1_not_7881_comb = ~p1_has_pos_inf__1_comb;
  assign p1_in0_r_sign__2_comb = p0_in0_r[31:31];
  assign p1_in0_i_sign__2_comb = p0_in0_i[31:31];

  // Registers for pipe stage 1:
  reg [7:0] p1_greater_exp_bexp;
  reg [7:0] p1_greater_exp_bexp__1;
  reg p1_greater_exp_sign;
  reg p1_greater_exp_sign__1;
  reg [27:0] p1_bit_slice_7808;
  reg [27:0] p1_bit_slice_7809;
  reg p1_bit_slice_7810;
  reg p1_bit_slice_7811;
  reg p1_ne_7814;
  reg p1_ne_7815;
  reg p1_nor_7860;
  reg p1_nor_7864;
  reg p1_is_result_nan__5;
  reg p1_is_operand_inf;
  reg p1_is_result_nan__6;
  reg p1_is_operand_inf__1;
  reg [22:0] p1_in0_r_fraction__6;
  reg [7:0] p1_in0_r_bexp__6;
  reg [22:0] p1_in0_i_fraction__6;
  reg [7:0] p1_in0_i_bexp__6;
  reg p1_fraction_is_zero;
  reg p1_fraction_is_zero__1;
  reg p1_not_7880;
  reg p1_not_7881;
  reg p1_in0_r_sign__2;
  reg p1_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p1_greater_exp_bexp <= p1_greater_exp_bexp_comb;
    p1_greater_exp_bexp__1 <= p1_greater_exp_bexp__1_comb;
    p1_greater_exp_sign <= p1_greater_exp_sign_comb;
    p1_greater_exp_sign__1 <= p1_greater_exp_sign__1_comb;
    p1_bit_slice_7808 <= p1_bit_slice_7808_comb;
    p1_bit_slice_7809 <= p1_bit_slice_7809_comb;
    p1_bit_slice_7810 <= p1_bit_slice_7810_comb;
    p1_bit_slice_7811 <= p1_bit_slice_7811_comb;
    p1_ne_7814 <= p1_ne_7814_comb;
    p1_ne_7815 <= p1_ne_7815_comb;
    p1_nor_7860 <= p1_nor_7860_comb;
    p1_nor_7864 <= p1_nor_7864_comb;
    p1_is_result_nan__5 <= p1_is_result_nan__5_comb;
    p1_is_operand_inf <= p1_is_operand_inf_comb;
    p1_is_result_nan__6 <= p1_is_result_nan__6_comb;
    p1_is_operand_inf__1 <= p1_is_operand_inf__1_comb;
    p1_in0_r_fraction__6 <= p1_in0_r_fraction__6_comb;
    p1_in0_r_bexp__6 <= p1_in0_r_bexp__6_comb;
    p1_in0_i_fraction__6 <= p1_in0_i_fraction__6_comb;
    p1_in0_i_bexp__6 <= p1_in0_i_bexp__6_comb;
    p1_fraction_is_zero <= p1_fraction_is_zero_comb;
    p1_fraction_is_zero__1 <= p1_fraction_is_zero__1_comb;
    p1_not_7880 <= p1_not_7880_comb;
    p1_not_7881 <= p1_not_7881_comb;
    p1_in0_r_sign__2 <= p1_in0_r_sign__2_comb;
    p1_in0_i_sign__2 <= p1_in0_i_sign__2_comb;
  end

  // ===== Pipe stage 2:
  wire [27:0] p2_abs_fraction_comb;
  wire [27:0] p2_abs_fraction__1_comb;
  wire [27:0] p2_reverse_7940_comb;
  wire [27:0] p2_reverse_7941_comb;
  wire [28:0] p2_one_hot_7942_comb;
  wire [28:0] p2_one_hot_7943_comb;
  wire [4:0] p2_encode_7944_comb;
  wire [4:0] p2_encode_7945_comb;
  wire p2_carry_bit_comb;
  wire p2_cancel_comb;
  wire p2_carry_bit__1_comb;
  wire p2_cancel__1_comb;
  wire [27:0] p2_leading_zeroes_comb;
  wire [27:0] p2_leading_zeroes__1_comb;
  wire [26:0] p2_carry_fraction_comb;
  wire [27:0] p2_add_7978_comb;
  wire [26:0] p2_carry_fraction__2_comb;
  wire [27:0] p2_add_7985_comb;
  wire [2:0] p2_concat_7986_comb;
  wire [26:0] p2_carry_fraction__1_comb;
  wire [26:0] p2_cancel_fraction_comb;
  wire [2:0] p2_concat_7989_comb;
  wire [26:0] p2_carry_fraction__3_comb;
  wire [26:0] p2_cancel_fraction__1_comb;
  wire [26:0] p2_shifted_fraction_comb;
  wire [26:0] p2_shifted_fraction__1_comb;
  wire [2:0] p2_normal_chunk_comb;
  wire [1:0] p2_half_way_chunk_comb;
  wire [2:0] p2_normal_chunk__1_comb;
  wire [1:0] p2_half_way_chunk__1_comb;
  wire [24:0] p2_add_8013_comb;
  wire [24:0] p2_add_8017_comb;
  wire p2_do_round_up__5_comb;
  wire p2_do_round_up__6_comb;
  wire [27:0] p2_rounded_fraction_comb;
  wire [27:0] p2_rounded_fraction__1_comb;
  wire p2_rounding_carry_comb;
  wire p2_rounding_carry__1_comb;
  wire [8:0] p2_add_8037_comb;
  wire [8:0] p2_add_8039_comb;
  wire [9:0] p2_add_8046_comb;
  wire [9:0] p2_add_8048_comb;
  wire [9:0] p2_wide_exponent_comb;
  wire [9:0] p2_wide_exponent__3_comb;
  wire [9:0] p2_wide_exponent__1_comb;
  wire [9:0] p2_wide_exponent__4_comb;
  wire [8:0] p2_wide_exponent__2_comb;
  wire [8:0] p2_wide_exponent__5_comb;
  wire [2:0] p2_add_8092_comb;
  wire [2:0] p2_add_8095_comb;
  wire [27:0] p2_shrl_8098_comb;
  wire p2_nor_8100_comb;
  wire [27:0] p2_shrl_8101_comb;
  wire p2_nor_8103_comb;
  wire [22:0] p2_result_fraction__13_comb;
  wire [22:0] p2_result_fraction__15_comb;
  wire [22:0] p2_result_fraction__14_comb;
  wire [22:0] p2_nan_fraction__14_comb;
  wire [7:0] p2_high_exp__36_comb;
  wire [22:0] p2_result_fraction__16_comb;
  wire [22:0] p2_nan_fraction__15_comb;
  wire [7:0] p2_high_exp__37_comb;
  wire [22:0] p2_result_fraction__17_comb;
  wire [7:0] p2_result_exponent__2_comb;
  wire [22:0] p2_result_fraction__18_comb;
  wire [7:0] p2_result_exponent__1_comb;
  wire [5:0] p2_add_8155_comb;
  wire p2_ugt_8157_comb;
  wire [5:0] p2_add_8166_comb;
  wire p2_ugt_8168_comb;
  wire p2_result_sign__9_comb;
  wire p2_result_sign__11_comb;
  wire [5:0] p2_add_8161_comb;
  wire [5:0] p2_add_8172_comb;
  wire [27:0] p2_wide_x__4_comb;
  wire [7:0] p2_greater_exp_bexp__2_comb;
  wire [27:0] p2_wide_x__6_comb;
  wire [7:0] p2_greater_exp_bexp__3_comb;
  wire [7:0] p2_high_exp__39_comb;
  wire p2_result_sign__10_comb;
  wire [7:0] p2_high_exp__41_comb;
  wire p2_result_sign__12_comb;
  wire [27:0] p2_wide_y__4_comb;
  wire [27:0] p2_wide_y__6_comb;
  wire [27:0] p2_wide_x__5_comb;
  wire [7:0] p2_sub_8193_comb;
  wire [27:0] p2_wide_x__7_comb;
  wire [7:0] p2_sub_8197_comb;
  wire [7:0] p2_high_exp__46_comb;
  wire p2_eq_8254_comb;
  wire p2_eq_8255_comb;
  wire [7:0] p2_high_exp__38_comb;
  wire p2_result_sign__13_comb;
  wire [7:0] p2_high_exp__47_comb;
  wire p2_eq_8260_comb;
  wire p2_eq_8261_comb;
  wire [7:0] p2_high_exp__40_comb;
  wire p2_result_sign__14_comb;
  wire [27:0] p2_wide_y__5_comb;
  wire [7:0] p2_sub_8195_comb;
  wire [27:0] p2_wide_y__7_comb;
  wire [7:0] p2_sub_8199_comb;
  wire [27:0] p2_dropped_x__2_comb;
  wire [27:0] p2_dropped_x__3_comb;
  wire p2_ne_8265_comb;
  wire p2_nand_8266_comb;
  wire p2_eq_8267_comb;
  wire p2_eq_8268_comb;
  wire p2_re__1_sign_comb;
  wire p2_ne_8270_comb;
  wire p2_nand_8271_comb;
  wire p2_eq_8272_comb;
  wire p2_eq_8273_comb;
  wire p2_im__1_sign_comb;
  wire [27:0] p2_dropped_y__2_comb;
  wire [27:0] p2_dropped_y__3_comb;
  wire p2_nor_8275_comb;
  wire p2_nor_8276_comb;
  wire p2_and_8277_comb;
  wire p2_nor_8278_comb;
  wire p2_nor_8280_comb;
  wire p2_nor_8281_comb;
  wire p2_and_8282_comb;
  wire p2_nor_8283_comb;
  wire [7:0] p2_shift_x__2_comb;
  wire p2_sticky_x__2_comb;
  wire [7:0] p2_shift_x__3_comb;
  wire p2_sticky_x__3_comb;
  wire p2_has_pos_inf__2_comb;
  wire p2_has_neg_inf__2_comb;
  wire p2_has_pos_inf__3_comb;
  wire p2_has_neg_inf__3_comb;
  wire p2_has_pos_inf__4_comb;
  wire p2_has_neg_inf__4_comb;
  wire p2_has_pos_inf__5_comb;
  wire p2_has_neg_inf__5_comb;
  wire [7:0] p2_shift_y__2_comb;
  wire p2_sticky_y__2_comb;
  wire [7:0] p2_shift_y__3_comb;
  wire p2_sticky_y__3_comb;
  wire [27:0] p2_shifted_x__2_comb;
  wire [27:0] p2_shifted_x__3_comb;
  wire p2_and_8287_comb;
  wire p2_and_8288_comb;
  wire p2_and_8292_comb;
  wire p2_and_8293_comb;
  wire p2_and_8298_comb;
  wire p2_and_8299_comb;
  wire p2_and_8302_comb;
  wire p2_and_8303_comb;
  wire [27:0] p2_shifted_y__2_comb;
  wire [27:0] p2_concat_8239_comb;
  wire [27:0] p2_shifted_y__3_comb;
  wire [27:0] p2_concat_8243_comb;
  wire [27:0] p2_addend_x__4_comb;
  wire [27:0] p2_addend_x__6_comb;
  wire p2_nor_8301_comb;
  wire p2_nor_8305_comb;
  wire p2_is_result_nan__7_comb;
  wire p2_is_operand_inf__2_comb;
  wire p2_not_8310_comb;
  wire p2_is_result_nan__8_comb;
  wire p2_is_operand_inf__3_comb;
  wire p2_not_8313_comb;
  wire p2_is_result_nan__9_comb;
  wire p2_not_8315_comb;
  wire p2_is_result_nan__10_comb;
  wire p2_not_8317_comb;
  assign p2_abs_fraction_comb = p1_bit_slice_7810 ? -p1_bit_slice_7808 : p1_bit_slice_7808;
  assign p2_abs_fraction__1_comb = p1_bit_slice_7811 ? -p1_bit_slice_7809 : p1_bit_slice_7809;
  assign p2_reverse_7940_comb = {p2_abs_fraction_comb[0], p2_abs_fraction_comb[1], p2_abs_fraction_comb[2], p2_abs_fraction_comb[3], p2_abs_fraction_comb[4], p2_abs_fraction_comb[5], p2_abs_fraction_comb[6], p2_abs_fraction_comb[7], p2_abs_fraction_comb[8], p2_abs_fraction_comb[9], p2_abs_fraction_comb[10], p2_abs_fraction_comb[11], p2_abs_fraction_comb[12], p2_abs_fraction_comb[13], p2_abs_fraction_comb[14], p2_abs_fraction_comb[15], p2_abs_fraction_comb[16], p2_abs_fraction_comb[17], p2_abs_fraction_comb[18], p2_abs_fraction_comb[19], p2_abs_fraction_comb[20], p2_abs_fraction_comb[21], p2_abs_fraction_comb[22], p2_abs_fraction_comb[23], p2_abs_fraction_comb[24], p2_abs_fraction_comb[25], p2_abs_fraction_comb[26], p2_abs_fraction_comb[27]};
  assign p2_reverse_7941_comb = {p2_abs_fraction__1_comb[0], p2_abs_fraction__1_comb[1], p2_abs_fraction__1_comb[2], p2_abs_fraction__1_comb[3], p2_abs_fraction__1_comb[4], p2_abs_fraction__1_comb[5], p2_abs_fraction__1_comb[6], p2_abs_fraction__1_comb[7], p2_abs_fraction__1_comb[8], p2_abs_fraction__1_comb[9], p2_abs_fraction__1_comb[10], p2_abs_fraction__1_comb[11], p2_abs_fraction__1_comb[12], p2_abs_fraction__1_comb[13], p2_abs_fraction__1_comb[14], p2_abs_fraction__1_comb[15], p2_abs_fraction__1_comb[16], p2_abs_fraction__1_comb[17], p2_abs_fraction__1_comb[18], p2_abs_fraction__1_comb[19], p2_abs_fraction__1_comb[20], p2_abs_fraction__1_comb[21], p2_abs_fraction__1_comb[22], p2_abs_fraction__1_comb[23], p2_abs_fraction__1_comb[24], p2_abs_fraction__1_comb[25], p2_abs_fraction__1_comb[26], p2_abs_fraction__1_comb[27]};
  assign p2_one_hot_7942_comb = {p2_reverse_7940_comb[27:0] == 28'h000_0000, p2_reverse_7940_comb[27] && p2_reverse_7940_comb[26:0] == 27'h000_0000, p2_reverse_7940_comb[26] && p2_reverse_7940_comb[25:0] == 26'h000_0000, p2_reverse_7940_comb[25] && p2_reverse_7940_comb[24:0] == 25'h000_0000, p2_reverse_7940_comb[24] && p2_reverse_7940_comb[23:0] == 24'h00_0000, p2_reverse_7940_comb[23] && p2_reverse_7940_comb[22:0] == 23'h00_0000, p2_reverse_7940_comb[22] && p2_reverse_7940_comb[21:0] == 22'h00_0000, p2_reverse_7940_comb[21] && p2_reverse_7940_comb[20:0] == 21'h00_0000, p2_reverse_7940_comb[20] && p2_reverse_7940_comb[19:0] == 20'h0_0000, p2_reverse_7940_comb[19] && p2_reverse_7940_comb[18:0] == 19'h0_0000, p2_reverse_7940_comb[18] && p2_reverse_7940_comb[17:0] == 18'h0_0000, p2_reverse_7940_comb[17] && p2_reverse_7940_comb[16:0] == 17'h0_0000, p2_reverse_7940_comb[16] && p2_reverse_7940_comb[15:0] == 16'h0000, p2_reverse_7940_comb[15] && p2_reverse_7940_comb[14:0] == 15'h0000, p2_reverse_7940_comb[14] && p2_reverse_7940_comb[13:0] == 14'h0000, p2_reverse_7940_comb[13] && p2_reverse_7940_comb[12:0] == 13'h0000, p2_reverse_7940_comb[12] && p2_reverse_7940_comb[11:0] == 12'h000, p2_reverse_7940_comb[11] && p2_reverse_7940_comb[10:0] == 11'h000, p2_reverse_7940_comb[10] && p2_reverse_7940_comb[9:0] == 10'h000, p2_reverse_7940_comb[9] && p2_reverse_7940_comb[8:0] == 9'h000, p2_reverse_7940_comb[8] && p2_reverse_7940_comb[7:0] == 8'h00, p2_reverse_7940_comb[7] && p2_reverse_7940_comb[6:0] == 7'h00, p2_reverse_7940_comb[6] && p2_reverse_7940_comb[5:0] == 6'h00, p2_reverse_7940_comb[5] && p2_reverse_7940_comb[4:0] == 5'h00, p2_reverse_7940_comb[4] && p2_reverse_7940_comb[3:0] == 4'h0, p2_reverse_7940_comb[3] && p2_reverse_7940_comb[2:0] == 3'h0, p2_reverse_7940_comb[2] && p2_reverse_7940_comb[1:0] == 2'h0, p2_reverse_7940_comb[1] && !p2_reverse_7940_comb[0], p2_reverse_7940_comb[0]};
  assign p2_one_hot_7943_comb = {p2_reverse_7941_comb[27:0] == 28'h000_0000, p2_reverse_7941_comb[27] && p2_reverse_7941_comb[26:0] == 27'h000_0000, p2_reverse_7941_comb[26] && p2_reverse_7941_comb[25:0] == 26'h000_0000, p2_reverse_7941_comb[25] && p2_reverse_7941_comb[24:0] == 25'h000_0000, p2_reverse_7941_comb[24] && p2_reverse_7941_comb[23:0] == 24'h00_0000, p2_reverse_7941_comb[23] && p2_reverse_7941_comb[22:0] == 23'h00_0000, p2_reverse_7941_comb[22] && p2_reverse_7941_comb[21:0] == 22'h00_0000, p2_reverse_7941_comb[21] && p2_reverse_7941_comb[20:0] == 21'h00_0000, p2_reverse_7941_comb[20] && p2_reverse_7941_comb[19:0] == 20'h0_0000, p2_reverse_7941_comb[19] && p2_reverse_7941_comb[18:0] == 19'h0_0000, p2_reverse_7941_comb[18] && p2_reverse_7941_comb[17:0] == 18'h0_0000, p2_reverse_7941_comb[17] && p2_reverse_7941_comb[16:0] == 17'h0_0000, p2_reverse_7941_comb[16] && p2_reverse_7941_comb[15:0] == 16'h0000, p2_reverse_7941_comb[15] && p2_reverse_7941_comb[14:0] == 15'h0000, p2_reverse_7941_comb[14] && p2_reverse_7941_comb[13:0] == 14'h0000, p2_reverse_7941_comb[13] && p2_reverse_7941_comb[12:0] == 13'h0000, p2_reverse_7941_comb[12] && p2_reverse_7941_comb[11:0] == 12'h000, p2_reverse_7941_comb[11] && p2_reverse_7941_comb[10:0] == 11'h000, p2_reverse_7941_comb[10] && p2_reverse_7941_comb[9:0] == 10'h000, p2_reverse_7941_comb[9] && p2_reverse_7941_comb[8:0] == 9'h000, p2_reverse_7941_comb[8] && p2_reverse_7941_comb[7:0] == 8'h00, p2_reverse_7941_comb[7] && p2_reverse_7941_comb[6:0] == 7'h00, p2_reverse_7941_comb[6] && p2_reverse_7941_comb[5:0] == 6'h00, p2_reverse_7941_comb[5] && p2_reverse_7941_comb[4:0] == 5'h00, p2_reverse_7941_comb[4] && p2_reverse_7941_comb[3:0] == 4'h0, p2_reverse_7941_comb[3] && p2_reverse_7941_comb[2:0] == 3'h0, p2_reverse_7941_comb[2] && p2_reverse_7941_comb[1:0] == 2'h0, p2_reverse_7941_comb[1] && !p2_reverse_7941_comb[0], p2_reverse_7941_comb[0]};
  assign p2_encode_7944_comb = {p2_one_hot_7942_comb[16] | p2_one_hot_7942_comb[17] | p2_one_hot_7942_comb[18] | p2_one_hot_7942_comb[19] | p2_one_hot_7942_comb[20] | p2_one_hot_7942_comb[21] | p2_one_hot_7942_comb[22] | p2_one_hot_7942_comb[23] | p2_one_hot_7942_comb[24] | p2_one_hot_7942_comb[25] | p2_one_hot_7942_comb[26] | p2_one_hot_7942_comb[27] | p2_one_hot_7942_comb[28], p2_one_hot_7942_comb[8] | p2_one_hot_7942_comb[9] | p2_one_hot_7942_comb[10] | p2_one_hot_7942_comb[11] | p2_one_hot_7942_comb[12] | p2_one_hot_7942_comb[13] | p2_one_hot_7942_comb[14] | p2_one_hot_7942_comb[15] | p2_one_hot_7942_comb[24] | p2_one_hot_7942_comb[25] | p2_one_hot_7942_comb[26] | p2_one_hot_7942_comb[27] | p2_one_hot_7942_comb[28], p2_one_hot_7942_comb[4] | p2_one_hot_7942_comb[5] | p2_one_hot_7942_comb[6] | p2_one_hot_7942_comb[7] | p2_one_hot_7942_comb[12] | p2_one_hot_7942_comb[13] | p2_one_hot_7942_comb[14] | p2_one_hot_7942_comb[15] | p2_one_hot_7942_comb[20] | p2_one_hot_7942_comb[21] | p2_one_hot_7942_comb[22] | p2_one_hot_7942_comb[23] | p2_one_hot_7942_comb[28], p2_one_hot_7942_comb[2] | p2_one_hot_7942_comb[3] | p2_one_hot_7942_comb[6] | p2_one_hot_7942_comb[7] | p2_one_hot_7942_comb[10] | p2_one_hot_7942_comb[11] | p2_one_hot_7942_comb[14] | p2_one_hot_7942_comb[15] | p2_one_hot_7942_comb[18] | p2_one_hot_7942_comb[19] | p2_one_hot_7942_comb[22] | p2_one_hot_7942_comb[23] | p2_one_hot_7942_comb[26] | p2_one_hot_7942_comb[27], p2_one_hot_7942_comb[1] | p2_one_hot_7942_comb[3] | p2_one_hot_7942_comb[5] | p2_one_hot_7942_comb[7] | p2_one_hot_7942_comb[9] | p2_one_hot_7942_comb[11] | p2_one_hot_7942_comb[13] | p2_one_hot_7942_comb[15] | p2_one_hot_7942_comb[17] | p2_one_hot_7942_comb[19] | p2_one_hot_7942_comb[21] | p2_one_hot_7942_comb[23] | p2_one_hot_7942_comb[25] | p2_one_hot_7942_comb[27]};
  assign p2_encode_7945_comb = {p2_one_hot_7943_comb[16] | p2_one_hot_7943_comb[17] | p2_one_hot_7943_comb[18] | p2_one_hot_7943_comb[19] | p2_one_hot_7943_comb[20] | p2_one_hot_7943_comb[21] | p2_one_hot_7943_comb[22] | p2_one_hot_7943_comb[23] | p2_one_hot_7943_comb[24] | p2_one_hot_7943_comb[25] | p2_one_hot_7943_comb[26] | p2_one_hot_7943_comb[27] | p2_one_hot_7943_comb[28], p2_one_hot_7943_comb[8] | p2_one_hot_7943_comb[9] | p2_one_hot_7943_comb[10] | p2_one_hot_7943_comb[11] | p2_one_hot_7943_comb[12] | p2_one_hot_7943_comb[13] | p2_one_hot_7943_comb[14] | p2_one_hot_7943_comb[15] | p2_one_hot_7943_comb[24] | p2_one_hot_7943_comb[25] | p2_one_hot_7943_comb[26] | p2_one_hot_7943_comb[27] | p2_one_hot_7943_comb[28], p2_one_hot_7943_comb[4] | p2_one_hot_7943_comb[5] | p2_one_hot_7943_comb[6] | p2_one_hot_7943_comb[7] | p2_one_hot_7943_comb[12] | p2_one_hot_7943_comb[13] | p2_one_hot_7943_comb[14] | p2_one_hot_7943_comb[15] | p2_one_hot_7943_comb[20] | p2_one_hot_7943_comb[21] | p2_one_hot_7943_comb[22] | p2_one_hot_7943_comb[23] | p2_one_hot_7943_comb[28], p2_one_hot_7943_comb[2] | p2_one_hot_7943_comb[3] | p2_one_hot_7943_comb[6] | p2_one_hot_7943_comb[7] | p2_one_hot_7943_comb[10] | p2_one_hot_7943_comb[11] | p2_one_hot_7943_comb[14] | p2_one_hot_7943_comb[15] | p2_one_hot_7943_comb[18] | p2_one_hot_7943_comb[19] | p2_one_hot_7943_comb[22] | p2_one_hot_7943_comb[23] | p2_one_hot_7943_comb[26] | p2_one_hot_7943_comb[27], p2_one_hot_7943_comb[1] | p2_one_hot_7943_comb[3] | p2_one_hot_7943_comb[5] | p2_one_hot_7943_comb[7] | p2_one_hot_7943_comb[9] | p2_one_hot_7943_comb[11] | p2_one_hot_7943_comb[13] | p2_one_hot_7943_comb[15] | p2_one_hot_7943_comb[17] | p2_one_hot_7943_comb[19] | p2_one_hot_7943_comb[21] | p2_one_hot_7943_comb[23] | p2_one_hot_7943_comb[25] | p2_one_hot_7943_comb[27]};
  assign p2_carry_bit_comb = p2_abs_fraction_comb[27];
  assign p2_cancel_comb = p2_encode_7944_comb[1] | p2_encode_7944_comb[2] | p2_encode_7944_comb[3] | p2_encode_7944_comb[4];
  assign p2_carry_bit__1_comb = p2_abs_fraction__1_comb[27];
  assign p2_cancel__1_comb = p2_encode_7945_comb[1] | p2_encode_7945_comb[2] | p2_encode_7945_comb[3] | p2_encode_7945_comb[4];
  assign p2_leading_zeroes_comb = {23'h00_0000, p2_encode_7944_comb};
  assign p2_leading_zeroes__1_comb = {23'h00_0000, p2_encode_7945_comb};
  assign p2_carry_fraction_comb = p2_abs_fraction_comb[27:1];
  assign p2_add_7978_comb = p2_leading_zeroes_comb + 28'hfff_ffff;
  assign p2_carry_fraction__2_comb = p2_abs_fraction__1_comb[27:1];
  assign p2_add_7985_comb = p2_leading_zeroes__1_comb + 28'hfff_ffff;
  assign p2_concat_7986_comb = {~p2_carry_bit_comb & ~p2_cancel_comb, ~p2_carry_bit_comb & p2_cancel_comb, p2_carry_bit_comb & ~p2_cancel_comb};
  assign p2_carry_fraction__1_comb = p2_carry_fraction_comb | {26'h000_0000, p2_abs_fraction_comb[0]};
  assign p2_cancel_fraction_comb = p2_add_7978_comb >= 28'h000_001b ? 27'h000_0000 : p2_abs_fraction_comb[26:0] << p2_add_7978_comb;
  assign p2_concat_7989_comb = {~p2_carry_bit__1_comb & ~p2_cancel__1_comb, ~p2_carry_bit__1_comb & p2_cancel__1_comb, p2_carry_bit__1_comb & ~p2_cancel__1_comb};
  assign p2_carry_fraction__3_comb = p2_carry_fraction__2_comb | {26'h000_0000, p2_abs_fraction__1_comb[0]};
  assign p2_cancel_fraction__1_comb = p2_add_7985_comb >= 28'h000_001b ? 27'h000_0000 : p2_abs_fraction__1_comb[26:0] << p2_add_7985_comb;
  assign p2_shifted_fraction_comb = p2_carry_fraction__1_comb & {27{p2_concat_7986_comb[0]}} | p2_cancel_fraction_comb & {27{p2_concat_7986_comb[1]}} | p2_abs_fraction_comb[26:0] & {27{p2_concat_7986_comb[2]}};
  assign p2_shifted_fraction__1_comb = p2_carry_fraction__3_comb & {27{p2_concat_7989_comb[0]}} | p2_cancel_fraction__1_comb & {27{p2_concat_7989_comb[1]}} | p2_abs_fraction__1_comb[26:0] & {27{p2_concat_7989_comb[2]}};
  assign p2_normal_chunk_comb = p2_shifted_fraction_comb[2:0];
  assign p2_half_way_chunk_comb = p2_shifted_fraction_comb[3:2];
  assign p2_normal_chunk__1_comb = p2_shifted_fraction__1_comb[2:0];
  assign p2_half_way_chunk__1_comb = p2_shifted_fraction__1_comb[3:2];
  assign p2_add_8013_comb = {1'h0, p2_shifted_fraction_comb[26:3]} + 25'h000_0001;
  assign p2_add_8017_comb = {1'h0, p2_shifted_fraction__1_comb[26:3]} + 25'h000_0001;
  assign p2_do_round_up__5_comb = p2_normal_chunk_comb > 3'h4 | p2_half_way_chunk_comb == 2'h3;
  assign p2_do_round_up__6_comb = p2_normal_chunk__1_comb > 3'h4 | p2_half_way_chunk__1_comb == 2'h3;
  assign p2_rounded_fraction_comb = p2_do_round_up__5_comb ? {p2_add_8013_comb, p2_normal_chunk_comb} : {1'h0, p2_shifted_fraction_comb};
  assign p2_rounded_fraction__1_comb = p2_do_round_up__6_comb ? {p2_add_8017_comb, p2_normal_chunk__1_comb} : {1'h0, p2_shifted_fraction__1_comb};
  assign p2_rounding_carry_comb = p2_rounded_fraction_comb[27];
  assign p2_rounding_carry__1_comb = p2_rounded_fraction__1_comb[27];
  assign p2_add_8037_comb = {1'h0, p1_greater_exp_bexp} + {8'h00, p2_rounding_carry_comb};
  assign p2_add_8039_comb = {1'h0, p1_greater_exp_bexp__1} + {8'h00, p2_rounding_carry__1_comb};
  assign p2_add_8046_comb = {1'h0, p2_add_8037_comb} + 10'h001;
  assign p2_add_8048_comb = {1'h0, p2_add_8039_comb} + 10'h001;
  assign p2_wide_exponent_comb = p2_add_8046_comb - {5'h00, p2_encode_7944_comb};
  assign p2_wide_exponent__3_comb = p2_add_8048_comb - {5'h00, p2_encode_7945_comb};
  assign p2_wide_exponent__1_comb = p2_wide_exponent_comb & {10{p1_ne_7814}};
  assign p2_wide_exponent__4_comb = p2_wide_exponent__3_comb & {10{p1_ne_7815}};
  assign p2_wide_exponent__2_comb = p2_wide_exponent__1_comb[8:0] & {9{~p2_wide_exponent__1_comb[9]}};
  assign p2_wide_exponent__5_comb = p2_wide_exponent__4_comb[8:0] & {9{~p2_wide_exponent__4_comb[9]}};
  assign p2_add_8092_comb = {2'h0, p2_rounding_carry_comb} + 3'h3;
  assign p2_add_8095_comb = {2'h0, p2_rounding_carry__1_comb} + 3'h3;
  assign p2_shrl_8098_comb = p2_rounded_fraction_comb >> p2_add_8092_comb;
  assign p2_nor_8100_comb = ~(p2_wide_exponent__2_comb[8] | p2_wide_exponent__2_comb[0] & p2_wide_exponent__2_comb[1] & p2_wide_exponent__2_comb[2] & p2_wide_exponent__2_comb[3] & p2_wide_exponent__2_comb[4] & p2_wide_exponent__2_comb[5] & p2_wide_exponent__2_comb[6] & p2_wide_exponent__2_comb[7]);
  assign p2_shrl_8101_comb = p2_rounded_fraction__1_comb >> p2_add_8095_comb;
  assign p2_nor_8103_comb = ~(p2_wide_exponent__5_comb[8] | p2_wide_exponent__5_comb[0] & p2_wide_exponent__5_comb[1] & p2_wide_exponent__5_comb[2] & p2_wide_exponent__5_comb[3] & p2_wide_exponent__5_comb[4] & p2_wide_exponent__5_comb[5] & p2_wide_exponent__5_comb[6] & p2_wide_exponent__5_comb[7]);
  assign p2_result_fraction__13_comb = p2_shrl_8098_comb[22:0];
  assign p2_result_fraction__15_comb = p2_shrl_8101_comb[22:0];
  assign p2_result_fraction__14_comb = p2_result_fraction__13_comb & {23{~(~(p2_wide_exponent__2_comb[1] | p2_wide_exponent__2_comb[2] | p2_wide_exponent__2_comb[3] | p2_wide_exponent__2_comb[4] | p2_wide_exponent__2_comb[5] | p2_wide_exponent__2_comb[6] | p2_wide_exponent__2_comb[7] | p2_wide_exponent__2_comb[8] | p2_wide_exponent__2_comb[0]))}} & {23{p2_nor_8100_comb}} & {23{p1_nor_7860}};
  assign p2_nan_fraction__14_comb = 23'h40_0000;
  assign p2_high_exp__36_comb = 8'hff;
  assign p2_result_fraction__16_comb = p2_result_fraction__15_comb & {23{~(~(p2_wide_exponent__5_comb[1] | p2_wide_exponent__5_comb[2] | p2_wide_exponent__5_comb[3] | p2_wide_exponent__5_comb[4] | p2_wide_exponent__5_comb[5] | p2_wide_exponent__5_comb[6] | p2_wide_exponent__5_comb[7] | p2_wide_exponent__5_comb[8] | p2_wide_exponent__5_comb[0]))}} & {23{p2_nor_8103_comb}} & {23{p1_nor_7864}};
  assign p2_nan_fraction__15_comb = 23'h40_0000;
  assign p2_high_exp__37_comb = 8'hff;
  assign p2_result_fraction__17_comb = p1_is_result_nan__5 ? p2_nan_fraction__14_comb : p2_result_fraction__14_comb;
  assign p2_result_exponent__2_comb = p1_is_result_nan__5 | p1_is_operand_inf | ~p2_nor_8100_comb ? p2_high_exp__36_comb : p2_wide_exponent__2_comb[7:0];
  assign p2_result_fraction__18_comb = p1_is_result_nan__6 ? p2_nan_fraction__15_comb : p2_result_fraction__16_comb;
  assign p2_result_exponent__1_comb = p1_is_result_nan__6 | p1_is_operand_inf__1 | ~p2_nor_8103_comb ? p2_high_exp__37_comb : p2_wide_exponent__5_comb[7:0];
  assign p2_add_8155_comb = p1_in0_r_bexp__6[7:2] + 6'h07;
  assign p2_ugt_8157_comb = p1_in0_r_bexp__6 > p2_result_exponent__2_comb;
  assign p2_add_8166_comb = p1_in0_i_bexp__6[7:2] + 6'h07;
  assign p2_ugt_8168_comb = p1_in0_i_bexp__6 > p2_result_exponent__1_comb;
  assign p2_result_sign__9_comb = ~(~p1_bit_slice_7810 | p1_greater_exp_sign) | ~(p1_bit_slice_7810 | p1_fraction_is_zero | ~p1_greater_exp_sign);
  assign p2_result_sign__11_comb = ~(~p1_bit_slice_7811 | p1_greater_exp_sign__1) | ~(p1_bit_slice_7811 | p1_fraction_is_zero__1 | ~p1_greater_exp_sign__1);
  assign p2_add_8161_comb = p2_result_exponent__2_comb[7:2] + 6'h07;
  assign p2_add_8172_comb = p2_result_exponent__1_comb[7:2] + 6'h07;
  assign p2_wide_x__4_comb = {{2'h0, p1_in0_r_fraction__6} | 25'h080_0000, 3'h0};
  assign p2_greater_exp_bexp__2_comb = p2_ugt_8157_comb ? p1_in0_r_bexp__6 : p2_result_exponent__2_comb;
  assign p2_wide_x__6_comb = {{2'h0, p1_in0_i_fraction__6} | 25'h080_0000, 3'h0};
  assign p2_greater_exp_bexp__3_comb = p2_ugt_8168_comb ? p1_in0_i_bexp__6 : p2_result_exponent__1_comb;
  assign p2_high_exp__39_comb = 8'hff;
  assign p2_result_sign__10_comb = p1_is_operand_inf ? p1_not_7880 : p2_result_sign__9_comb;
  assign p2_high_exp__41_comb = 8'hff;
  assign p2_result_sign__12_comb = p1_is_operand_inf__1 ? p1_not_7881 : p2_result_sign__11_comb;
  assign p2_wide_y__4_comb = {{2'h0, p2_result_fraction__17_comb} | 25'h080_0000, 3'h0};
  assign p2_wide_y__6_comb = {{2'h0, p2_result_fraction__18_comb} | 25'h080_0000, 3'h0};
  assign p2_wide_x__5_comb = p2_wide_x__4_comb & {28{p1_in0_r_bexp__6 != 8'h00}};
  assign p2_sub_8193_comb = {p2_add_8155_comb, p1_in0_r_bexp__6[1:0]} - p2_greater_exp_bexp__2_comb;
  assign p2_wide_x__7_comb = p2_wide_x__6_comb & {28{p1_in0_i_bexp__6 != 8'h00}};
  assign p2_sub_8197_comb = {p2_add_8166_comb, p1_in0_i_bexp__6[1:0]} - p2_greater_exp_bexp__3_comb;
  assign p2_high_exp__46_comb = 8'hff;
  assign p2_eq_8254_comb = p2_result_exponent__2_comb == p2_high_exp__39_comb;
  assign p2_eq_8255_comb = p2_result_fraction__17_comb == 23'h00_0000;
  assign p2_high_exp__38_comb = 8'hff;
  assign p2_result_sign__13_comb = ~p1_is_result_nan__5 & p2_result_sign__10_comb;
  assign p2_high_exp__47_comb = 8'hff;
  assign p2_eq_8260_comb = p2_result_exponent__1_comb == p2_high_exp__41_comb;
  assign p2_eq_8261_comb = p2_result_fraction__18_comb == 23'h00_0000;
  assign p2_high_exp__40_comb = 8'hff;
  assign p2_result_sign__14_comb = ~p1_is_result_nan__6 & p2_result_sign__12_comb;
  assign p2_wide_y__5_comb = p2_wide_y__4_comb & {28{p2_result_exponent__2_comb != 8'h00}};
  assign p2_sub_8195_comb = {p2_add_8161_comb, p2_result_exponent__2_comb[1:0]} - p2_greater_exp_bexp__2_comb;
  assign p2_wide_y__7_comb = p2_wide_y__6_comb & {28{p2_result_exponent__1_comb != 8'h00}};
  assign p2_sub_8199_comb = {p2_add_8172_comb, p2_result_exponent__1_comb[1:0]} - p2_greater_exp_bexp__3_comb;
  assign p2_dropped_x__2_comb = p2_sub_8193_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__5_comb << p2_sub_8193_comb;
  assign p2_dropped_x__3_comb = p2_sub_8197_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__7_comb << p2_sub_8197_comb;
  assign p2_ne_8265_comb = p1_in0_r_fraction__6 != 23'h00_0000;
  assign p2_nand_8266_comb = ~(p2_eq_8254_comb & p2_eq_8255_comb);
  assign p2_eq_8267_comb = p1_in0_r_bexp__6 == p2_high_exp__38_comb;
  assign p2_eq_8268_comb = p1_in0_r_fraction__6 == 23'h00_0000;
  assign p2_re__1_sign_comb = ~p2_result_sign__13_comb;
  assign p2_ne_8270_comb = p1_in0_i_fraction__6 != 23'h00_0000;
  assign p2_nand_8271_comb = ~(p2_eq_8260_comb & p2_eq_8261_comb);
  assign p2_eq_8272_comb = p1_in0_i_bexp__6 == p2_high_exp__40_comb;
  assign p2_eq_8273_comb = p1_in0_i_fraction__6 == 23'h00_0000;
  assign p2_im__1_sign_comb = ~p2_result_sign__14_comb;
  assign p2_dropped_y__2_comb = p2_sub_8195_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__5_comb << p2_sub_8195_comb;
  assign p2_dropped_y__3_comb = p2_sub_8199_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__7_comb << p2_sub_8199_comb;
  assign p2_nor_8275_comb = ~(p1_in0_r_bexp__6 != p2_high_exp__46_comb | p2_ne_8265_comb | p1_in0_r_sign__2);
  assign p2_nor_8276_comb = ~(p2_nand_8266_comb | p2_result_sign__13_comb);
  assign p2_and_8277_comb = p2_eq_8267_comb & p2_eq_8268_comb & p1_in0_r_sign__2;
  assign p2_nor_8278_comb = ~(p2_nand_8266_comb | p2_re__1_sign_comb);
  assign p2_nor_8280_comb = ~(p1_in0_i_bexp__6 != p2_high_exp__47_comb | p2_ne_8270_comb | p1_in0_i_sign__2);
  assign p2_nor_8281_comb = ~(p2_nand_8271_comb | p2_result_sign__14_comb);
  assign p2_and_8282_comb = p2_eq_8272_comb & p2_eq_8273_comb & p1_in0_i_sign__2;
  assign p2_nor_8283_comb = ~(p2_nand_8271_comb | p2_im__1_sign_comb);
  assign p2_shift_x__2_comb = p2_greater_exp_bexp__2_comb - p1_in0_r_bexp__6;
  assign p2_sticky_x__2_comb = p2_dropped_x__2_comb[27:3] != 25'h000_0000;
  assign p2_shift_x__3_comb = p2_greater_exp_bexp__3_comb - p1_in0_i_bexp__6;
  assign p2_sticky_x__3_comb = p2_dropped_x__3_comb[27:3] != 25'h000_0000;
  assign p2_has_pos_inf__2_comb = p2_nor_8275_comb | p2_nor_8276_comb;
  assign p2_has_neg_inf__2_comb = p2_and_8277_comb | p2_nor_8278_comb;
  assign p2_has_pos_inf__3_comb = p2_nor_8280_comb | p2_nor_8281_comb;
  assign p2_has_neg_inf__3_comb = p2_and_8282_comb | p2_nor_8283_comb;
  assign p2_has_pos_inf__4_comb = p2_nor_8275_comb | p2_nor_8278_comb;
  assign p2_has_neg_inf__4_comb = p2_and_8277_comb | p2_nor_8276_comb;
  assign p2_has_pos_inf__5_comb = p2_nor_8280_comb | p2_nor_8283_comb;
  assign p2_has_neg_inf__5_comb = p2_and_8282_comb | p2_nor_8281_comb;
  assign p2_shift_y__2_comb = p2_greater_exp_bexp__2_comb - p2_result_exponent__2_comb;
  assign p2_sticky_y__2_comb = p2_dropped_y__2_comb[27:3] != 25'h000_0000;
  assign p2_shift_y__3_comb = p2_greater_exp_bexp__3_comb - p2_result_exponent__1_comb;
  assign p2_sticky_y__3_comb = p2_dropped_y__3_comb[27:3] != 25'h000_0000;
  assign p2_shifted_x__2_comb = p2_shift_x__2_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__5_comb >> p2_shift_x__2_comb;
  assign p2_shifted_x__3_comb = p2_shift_x__3_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__7_comb >> p2_shift_x__3_comb;
  assign p2_and_8287_comb = p2_eq_8267_comb & p2_eq_8268_comb;
  assign p2_and_8288_comb = p2_eq_8254_comb & p2_eq_8255_comb;
  assign p2_and_8292_comb = p2_eq_8272_comb & p2_eq_8273_comb;
  assign p2_and_8293_comb = p2_eq_8260_comb & p2_eq_8261_comb;
  assign p2_and_8298_comb = p2_eq_8267_comb & p2_ne_8265_comb;
  assign p2_and_8299_comb = p2_eq_8254_comb & p2_result_fraction__17_comb != 23'h00_0000;
  assign p2_and_8302_comb = p2_eq_8272_comb & p2_ne_8270_comb;
  assign p2_and_8303_comb = p2_eq_8260_comb & p2_result_fraction__18_comb != 23'h00_0000;
  assign p2_shifted_y__2_comb = p2_shift_y__2_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__5_comb >> p2_shift_y__2_comb;
  assign p2_concat_8239_comb = {27'h000_0000, p2_sticky_y__2_comb};
  assign p2_shifted_y__3_comb = p2_shift_y__3_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__7_comb >> p2_shift_y__3_comb;
  assign p2_concat_8243_comb = {27'h000_0000, p2_sticky_y__3_comb};
  assign p2_addend_x__4_comb = p2_shifted_x__2_comb | {27'h000_0000, p2_sticky_x__2_comb};
  assign p2_addend_x__6_comb = p2_shifted_x__3_comb | {27'h000_0000, p2_sticky_x__3_comb};
  assign p2_nor_8301_comb = ~(p2_and_8287_comb | p2_and_8288_comb);
  assign p2_nor_8305_comb = ~(p2_and_8292_comb | p2_and_8293_comb);
  assign p2_is_result_nan__7_comb = p2_and_8298_comb | p2_and_8299_comb | p2_has_pos_inf__2_comb & p2_has_neg_inf__2_comb;
  assign p2_is_operand_inf__2_comb = p2_and_8287_comb | p2_and_8288_comb;
  assign p2_not_8310_comb = ~p2_has_pos_inf__2_comb;
  assign p2_is_result_nan__8_comb = p2_and_8302_comb | p2_and_8303_comb | p2_has_pos_inf__3_comb & p2_has_neg_inf__3_comb;
  assign p2_is_operand_inf__3_comb = p2_and_8292_comb | p2_and_8293_comb;
  assign p2_not_8313_comb = ~p2_has_pos_inf__3_comb;
  assign p2_is_result_nan__9_comb = p2_and_8298_comb | p2_and_8299_comb | p2_has_pos_inf__4_comb & p2_has_neg_inf__4_comb;
  assign p2_not_8315_comb = ~p2_has_pos_inf__4_comb;
  assign p2_is_result_nan__10_comb = p2_and_8302_comb | p2_and_8303_comb | p2_has_pos_inf__5_comb & p2_has_neg_inf__5_comb;
  assign p2_not_8317_comb = ~p2_has_pos_inf__5_comb;

  // Registers for pipe stage 2:
  reg p2_ugt_8157;
  reg p2_ugt_8168;
  reg [7:0] p2_greater_exp_bexp__2;
  reg [7:0] p2_greater_exp_bexp__3;
  reg p2_result_sign__13;
  reg p2_result_sign__14;
  reg p2_in0_r_sign__2;
  reg [27:0] p2_shifted_y__2;
  reg [27:0] p2_concat_8239;
  reg p2_in0_i_sign__2;
  reg [27:0] p2_shifted_y__3;
  reg [27:0] p2_concat_8243;
  reg p2_re__1_sign;
  reg p2_im__1_sign;
  reg [27:0] p2_addend_x__4;
  reg [27:0] p2_addend_x__6;
  reg p2_nor_8301;
  reg p2_nor_8305;
  reg p2_is_result_nan__7;
  reg p2_is_operand_inf__2;
  reg p2_not_8310;
  reg p2_is_result_nan__8;
  reg p2_is_operand_inf__3;
  reg p2_not_8313;
  reg p2_is_result_nan__9;
  reg p2_not_8315;
  reg p2_is_result_nan__10;
  reg p2_not_8317;
  always_ff @ (posedge clk) begin
    p2_ugt_8157 <= p2_ugt_8157_comb;
    p2_ugt_8168 <= p2_ugt_8168_comb;
    p2_greater_exp_bexp__2 <= p2_greater_exp_bexp__2_comb;
    p2_greater_exp_bexp__3 <= p2_greater_exp_bexp__3_comb;
    p2_result_sign__13 <= p2_result_sign__13_comb;
    p2_result_sign__14 <= p2_result_sign__14_comb;
    p2_in0_r_sign__2 <= p1_in0_r_sign__2;
    p2_shifted_y__2 <= p2_shifted_y__2_comb;
    p2_concat_8239 <= p2_concat_8239_comb;
    p2_in0_i_sign__2 <= p1_in0_i_sign__2;
    p2_shifted_y__3 <= p2_shifted_y__3_comb;
    p2_concat_8243 <= p2_concat_8243_comb;
    p2_re__1_sign <= p2_re__1_sign_comb;
    p2_im__1_sign <= p2_im__1_sign_comb;
    p2_addend_x__4 <= p2_addend_x__4_comb;
    p2_addend_x__6 <= p2_addend_x__6_comb;
    p2_nor_8301 <= p2_nor_8301_comb;
    p2_nor_8305 <= p2_nor_8305_comb;
    p2_is_result_nan__7 <= p2_is_result_nan__7_comb;
    p2_is_operand_inf__2 <= p2_is_operand_inf__2_comb;
    p2_not_8310 <= p2_not_8310_comb;
    p2_is_result_nan__8 <= p2_is_result_nan__8_comb;
    p2_is_operand_inf__3 <= p2_is_operand_inf__3_comb;
    p2_not_8313 <= p2_not_8313_comb;
    p2_is_result_nan__9 <= p2_is_result_nan__9_comb;
    p2_not_8315 <= p2_not_8315_comb;
    p2_is_result_nan__10 <= p2_is_result_nan__10_comb;
    p2_not_8317 <= p2_not_8317_comb;
  end

  // ===== Pipe stage 3:
  wire p3_greater_exp_sign__2_comb;
  wire [27:0] p3_addend_y__4_comb;
  wire p3_greater_exp_sign__3_comb;
  wire [27:0] p3_addend_y__6_comb;
  wire p3_greater_exp_sign__4_comb;
  wire p3_greater_exp_sign__5_comb;
  wire [27:0] p3_addend_x__5_comb;
  wire [27:0] p3_addend_y__5_comb;
  wire [27:0] p3_addend_x__7_comb;
  wire [27:0] p3_addend_y__7_comb;
  wire [27:0] p3_addend_x__9_comb;
  wire [27:0] p3_addend_y__9_comb;
  wire [27:0] p3_addend_x__11_comb;
  wire [27:0] p3_addend_y__11_comb;
  wire [28:0] p3_fraction__35_comb;
  wire [28:0] p3_fraction__36_comb;
  wire [28:0] p3_fraction__37_comb;
  wire [28:0] p3_fraction__38_comb;
  wire [27:0] p3_abs_fraction__2_comb;
  wire [27:0] p3_abs_fraction__3_comb;
  wire [27:0] p3_abs_fraction__4_comb;
  wire [27:0] p3_abs_fraction__5_comb;
  wire [27:0] p3_reverse_8428_comb;
  wire [27:0] p3_reverse_8429_comb;
  wire [27:0] p3_reverse_8430_comb;
  wire [27:0] p3_reverse_8431_comb;
  wire [28:0] p3_one_hot_8432_comb;
  wire [28:0] p3_one_hot_8433_comb;
  wire [28:0] p3_one_hot_8434_comb;
  wire [28:0] p3_one_hot_8435_comb;
  wire [4:0] p3_encode_8436_comb;
  wire [4:0] p3_encode_8437_comb;
  wire [4:0] p3_encode_8438_comb;
  wire [4:0] p3_encode_8439_comb;
  wire p3_carry_bit__2_comb;
  wire p3_cancel__2_comb;
  wire p3_carry_bit__3_comb;
  wire p3_cancel__3_comb;
  wire p3_carry_bit__4_comb;
  wire p3_cancel__4_comb;
  wire p3_carry_bit__5_comb;
  wire p3_cancel__5_comb;
  wire [27:0] p3_leading_zeroes__2_comb;
  wire [27:0] p3_leading_zeroes__3_comb;
  wire [27:0] p3_leading_zeroes__4_comb;
  wire [27:0] p3_leading_zeroes__5_comb;
  wire [26:0] p3_carry_fraction__4_comb;
  wire [27:0] p3_add_8498_comb;
  wire [26:0] p3_carry_fraction__6_comb;
  wire [27:0] p3_add_8505_comb;
  wire [26:0] p3_carry_fraction__8_comb;
  wire [27:0] p3_add_8512_comb;
  wire [26:0] p3_carry_fraction__10_comb;
  wire [27:0] p3_add_8519_comb;
  wire [2:0] p3_concat_8520_comb;
  wire [26:0] p3_carry_fraction__5_comb;
  wire [26:0] p3_cancel_fraction__2_comb;
  wire [2:0] p3_concat_8523_comb;
  wire [26:0] p3_carry_fraction__7_comb;
  wire [26:0] p3_cancel_fraction__3_comb;
  wire [2:0] p3_concat_8526_comb;
  wire [26:0] p3_carry_fraction__9_comb;
  wire [26:0] p3_cancel_fraction__4_comb;
  wire [2:0] p3_concat_8529_comb;
  wire [26:0] p3_carry_fraction__11_comb;
  wire [26:0] p3_cancel_fraction__5_comb;
  wire [26:0] p3_shifted_fraction__2_comb;
  wire [26:0] p3_shifted_fraction__3_comb;
  wire [26:0] p3_shifted_fraction__4_comb;
  wire [26:0] p3_shifted_fraction__5_comb;
  wire [2:0] p3_normal_chunk__2_comb;
  wire [1:0] p3_half_way_chunk__2_comb;
  wire [2:0] p3_normal_chunk__3_comb;
  wire [1:0] p3_half_way_chunk__3_comb;
  wire [2:0] p3_normal_chunk__4_comb;
  wire [1:0] p3_half_way_chunk__4_comb;
  wire [2:0] p3_normal_chunk__5_comb;
  wire [1:0] p3_half_way_chunk__5_comb;
  wire [24:0] p3_add_8571_comb;
  wire [24:0] p3_add_8575_comb;
  wire [24:0] p3_add_8579_comb;
  wire [24:0] p3_add_8583_comb;
  wire p3_do_round_up__7_comb;
  wire p3_do_round_up__8_comb;
  wire p3_do_round_up__9_comb;
  wire p3_do_round_up__10_comb;
  wire [27:0] p3_rounded_fraction__2_comb;
  wire [27:0] p3_rounded_fraction__3_comb;
  wire [27:0] p3_rounded_fraction__4_comb;
  wire [27:0] p3_rounded_fraction__5_comb;
  wire p3_rounding_carry__2_comb;
  wire p3_rounding_carry__3_comb;
  wire p3_rounding_carry__4_comb;
  wire p3_rounding_carry__5_comb;
  wire [8:0] p3_concat_8610_comb;
  wire [8:0] p3_concat_8612_comb;
  wire [8:0] p3_add_8617_comb;
  wire [8:0] p3_add_8619_comb;
  wire [8:0] p3_add_8621_comb;
  wire [8:0] p3_add_8623_comb;
  wire [9:0] p3_add_8640_comb;
  wire [9:0] p3_add_8643_comb;
  wire [9:0] p3_add_8646_comb;
  wire [9:0] p3_add_8649_comb;
  wire [9:0] p3_wide_exponent__6_comb;
  wire [9:0] p3_wide_exponent__9_comb;
  wire [9:0] p3_wide_exponent__12_comb;
  wire [9:0] p3_wide_exponent__15_comb;
  wire [9:0] p3_wide_exponent__7_comb;
  wire [9:0] p3_wide_exponent__10_comb;
  wire [9:0] p3_wide_exponent__13_comb;
  wire [9:0] p3_wide_exponent__16_comb;
  wire [8:0] p3_wide_exponent__8_comb;
  wire [8:0] p3_wide_exponent__11_comb;
  wire [8:0] p3_wide_exponent__14_comb;
  wire [8:0] p3_wide_exponent__17_comb;
  wire p3_fraction_is_zero__2_comb;
  wire [2:0] p3_add_8744_comb;
  wire p3_fraction_is_zero__3_comb;
  wire [2:0] p3_add_8750_comb;
  wire p3_fraction_is_zero__4_comb;
  wire [2:0] p3_add_8756_comb;
  wire p3_fraction_is_zero__5_comb;
  wire [2:0] p3_add_8762_comb;
  wire p3_nor_8766_comb;
  wire [27:0] p3_shrl_8767_comb;
  wire p3_nor_8771_comb;
  wire [27:0] p3_shrl_8772_comb;
  wire p3_nor_8776_comb;
  wire [27:0] p3_shrl_8777_comb;
  wire p3_nor_8781_comb;
  wire [27:0] p3_shrl_8782_comb;
  wire p3_result_sign__15_comb;
  wire [22:0] p3_result_fraction__19_comb;
  wire [22:0] p3_sign_ext_8789_comb;
  wire p3_result_sign__17_comb;
  wire [22:0] p3_result_fraction__21_comb;
  wire [22:0] p3_sign_ext_8795_comb;
  wire p3_result_sign__20_comb;
  wire [22:0] p3_result_fraction__24_comb;
  wire p3_result_sign__23_comb;
  wire [22:0] p3_result_fraction__27_comb;
  wire p3_result_sign__16_comb;
  wire [7:0] p3_high_exp__42_comb;
  wire [22:0] p3_result_fraction__20_comb;
  wire [22:0] p3_nan_fraction__16_comb;
  wire p3_result_sign__18_comb;
  wire [7:0] p3_high_exp__43_comb;
  wire [22:0] p3_result_fraction__22_comb;
  wire [22:0] p3_nan_fraction__17_comb;
  wire p3_result_sign__21_comb;
  wire [7:0] p3_high_exp__44_comb;
  wire [22:0] p3_result_fraction__25_comb;
  wire [22:0] p3_nan_fraction__18_comb;
  wire p3_result_sign__24_comb;
  wire [7:0] p3_high_exp__45_comb;
  wire [22:0] p3_result_fraction__28_comb;
  wire [22:0] p3_nan_fraction__19_comb;
  wire p3_result_sign__19_comb;
  wire [7:0] p3_result_exponent__3_comb;
  wire [22:0] p3_result_fraction__23_comb;
  wire p3_result_sign__22_comb;
  wire [7:0] p3_result_exponent__4_comb;
  wire [22:0] p3_result_fraction__26_comb;
  wire p3_result_sign__25_comb;
  wire [7:0] p3_result_exponent__5_comb;
  wire [22:0] p3_result_fraction__29_comb;
  wire p3_result_sign__26_comb;
  wire [7:0] p3_result_exponent__6_comb;
  wire [22:0] p3_result_fraction__30_comb;
  wire [31:0] p3_out0_r_comb;
  wire [31:0] p3_out0_i_comb;
  wire [31:0] p3_out1_r_comb;
  wire [31:0] p3_out1_i_comb;
  wire [127:0] p3_tuple_8850_comb;
  assign p3_greater_exp_sign__2_comb = p2_ugt_8157 ? p2_in0_r_sign__2 : p2_result_sign__13;
  assign p3_addend_y__4_comb = p2_shifted_y__2 | p2_concat_8239;
  assign p3_greater_exp_sign__3_comb = p2_ugt_8168 ? p2_in0_i_sign__2 : p2_result_sign__14;
  assign p3_addend_y__6_comb = p2_shifted_y__3 | p2_concat_8243;
  assign p3_greater_exp_sign__4_comb = p2_ugt_8157 ? p2_in0_r_sign__2 : p2_re__1_sign;
  assign p3_greater_exp_sign__5_comb = p2_ugt_8168 ? p2_in0_i_sign__2 : p2_im__1_sign;
  assign p3_addend_x__5_comb = p2_in0_r_sign__2 ^ p3_greater_exp_sign__2_comb ? -p2_addend_x__4 : p2_addend_x__4;
  assign p3_addend_y__5_comb = p2_result_sign__13 ^ p3_greater_exp_sign__2_comb ? -p3_addend_y__4_comb : p3_addend_y__4_comb;
  assign p3_addend_x__7_comb = p2_in0_i_sign__2 ^ p3_greater_exp_sign__3_comb ? -p2_addend_x__6 : p2_addend_x__6;
  assign p3_addend_y__7_comb = p2_result_sign__14 ^ p3_greater_exp_sign__3_comb ? -p3_addend_y__6_comb : p3_addend_y__6_comb;
  assign p3_addend_x__9_comb = p2_in0_r_sign__2 ^ p3_greater_exp_sign__4_comb ? -p2_addend_x__4 : p2_addend_x__4;
  assign p3_addend_y__9_comb = p2_re__1_sign ^ p3_greater_exp_sign__4_comb ? -p3_addend_y__4_comb : p3_addend_y__4_comb;
  assign p3_addend_x__11_comb = p2_in0_i_sign__2 ^ p3_greater_exp_sign__5_comb ? -p2_addend_x__6 : p2_addend_x__6;
  assign p3_addend_y__11_comb = p2_im__1_sign ^ p3_greater_exp_sign__5_comb ? -p3_addend_y__6_comb : p3_addend_y__6_comb;
  assign p3_fraction__35_comb = {{1{p3_addend_x__5_comb[27]}}, p3_addend_x__5_comb} + {{1{p3_addend_y__5_comb[27]}}, p3_addend_y__5_comb};
  assign p3_fraction__36_comb = {{1{p3_addend_x__7_comb[27]}}, p3_addend_x__7_comb} + {{1{p3_addend_y__7_comb[27]}}, p3_addend_y__7_comb};
  assign p3_fraction__37_comb = {{1{p3_addend_x__9_comb[27]}}, p3_addend_x__9_comb} + {{1{p3_addend_y__9_comb[27]}}, p3_addend_y__9_comb};
  assign p3_fraction__38_comb = {{1{p3_addend_x__11_comb[27]}}, p3_addend_x__11_comb} + {{1{p3_addend_y__11_comb[27]}}, p3_addend_y__11_comb};
  assign p3_abs_fraction__2_comb = p3_fraction__35_comb[28] ? -p3_fraction__35_comb[27:0] : p3_fraction__35_comb[27:0];
  assign p3_abs_fraction__3_comb = p3_fraction__36_comb[28] ? -p3_fraction__36_comb[27:0] : p3_fraction__36_comb[27:0];
  assign p3_abs_fraction__4_comb = p3_fraction__37_comb[28] ? -p3_fraction__37_comb[27:0] : p3_fraction__37_comb[27:0];
  assign p3_abs_fraction__5_comb = p3_fraction__38_comb[28] ? -p3_fraction__38_comb[27:0] : p3_fraction__38_comb[27:0];
  assign p3_reverse_8428_comb = {p3_abs_fraction__2_comb[0], p3_abs_fraction__2_comb[1], p3_abs_fraction__2_comb[2], p3_abs_fraction__2_comb[3], p3_abs_fraction__2_comb[4], p3_abs_fraction__2_comb[5], p3_abs_fraction__2_comb[6], p3_abs_fraction__2_comb[7], p3_abs_fraction__2_comb[8], p3_abs_fraction__2_comb[9], p3_abs_fraction__2_comb[10], p3_abs_fraction__2_comb[11], p3_abs_fraction__2_comb[12], p3_abs_fraction__2_comb[13], p3_abs_fraction__2_comb[14], p3_abs_fraction__2_comb[15], p3_abs_fraction__2_comb[16], p3_abs_fraction__2_comb[17], p3_abs_fraction__2_comb[18], p3_abs_fraction__2_comb[19], p3_abs_fraction__2_comb[20], p3_abs_fraction__2_comb[21], p3_abs_fraction__2_comb[22], p3_abs_fraction__2_comb[23], p3_abs_fraction__2_comb[24], p3_abs_fraction__2_comb[25], p3_abs_fraction__2_comb[26], p3_abs_fraction__2_comb[27]};
  assign p3_reverse_8429_comb = {p3_abs_fraction__3_comb[0], p3_abs_fraction__3_comb[1], p3_abs_fraction__3_comb[2], p3_abs_fraction__3_comb[3], p3_abs_fraction__3_comb[4], p3_abs_fraction__3_comb[5], p3_abs_fraction__3_comb[6], p3_abs_fraction__3_comb[7], p3_abs_fraction__3_comb[8], p3_abs_fraction__3_comb[9], p3_abs_fraction__3_comb[10], p3_abs_fraction__3_comb[11], p3_abs_fraction__3_comb[12], p3_abs_fraction__3_comb[13], p3_abs_fraction__3_comb[14], p3_abs_fraction__3_comb[15], p3_abs_fraction__3_comb[16], p3_abs_fraction__3_comb[17], p3_abs_fraction__3_comb[18], p3_abs_fraction__3_comb[19], p3_abs_fraction__3_comb[20], p3_abs_fraction__3_comb[21], p3_abs_fraction__3_comb[22], p3_abs_fraction__3_comb[23], p3_abs_fraction__3_comb[24], p3_abs_fraction__3_comb[25], p3_abs_fraction__3_comb[26], p3_abs_fraction__3_comb[27]};
  assign p3_reverse_8430_comb = {p3_abs_fraction__4_comb[0], p3_abs_fraction__4_comb[1], p3_abs_fraction__4_comb[2], p3_abs_fraction__4_comb[3], p3_abs_fraction__4_comb[4], p3_abs_fraction__4_comb[5], p3_abs_fraction__4_comb[6], p3_abs_fraction__4_comb[7], p3_abs_fraction__4_comb[8], p3_abs_fraction__4_comb[9], p3_abs_fraction__4_comb[10], p3_abs_fraction__4_comb[11], p3_abs_fraction__4_comb[12], p3_abs_fraction__4_comb[13], p3_abs_fraction__4_comb[14], p3_abs_fraction__4_comb[15], p3_abs_fraction__4_comb[16], p3_abs_fraction__4_comb[17], p3_abs_fraction__4_comb[18], p3_abs_fraction__4_comb[19], p3_abs_fraction__4_comb[20], p3_abs_fraction__4_comb[21], p3_abs_fraction__4_comb[22], p3_abs_fraction__4_comb[23], p3_abs_fraction__4_comb[24], p3_abs_fraction__4_comb[25], p3_abs_fraction__4_comb[26], p3_abs_fraction__4_comb[27]};
  assign p3_reverse_8431_comb = {p3_abs_fraction__5_comb[0], p3_abs_fraction__5_comb[1], p3_abs_fraction__5_comb[2], p3_abs_fraction__5_comb[3], p3_abs_fraction__5_comb[4], p3_abs_fraction__5_comb[5], p3_abs_fraction__5_comb[6], p3_abs_fraction__5_comb[7], p3_abs_fraction__5_comb[8], p3_abs_fraction__5_comb[9], p3_abs_fraction__5_comb[10], p3_abs_fraction__5_comb[11], p3_abs_fraction__5_comb[12], p3_abs_fraction__5_comb[13], p3_abs_fraction__5_comb[14], p3_abs_fraction__5_comb[15], p3_abs_fraction__5_comb[16], p3_abs_fraction__5_comb[17], p3_abs_fraction__5_comb[18], p3_abs_fraction__5_comb[19], p3_abs_fraction__5_comb[20], p3_abs_fraction__5_comb[21], p3_abs_fraction__5_comb[22], p3_abs_fraction__5_comb[23], p3_abs_fraction__5_comb[24], p3_abs_fraction__5_comb[25], p3_abs_fraction__5_comb[26], p3_abs_fraction__5_comb[27]};
  assign p3_one_hot_8432_comb = {p3_reverse_8428_comb[27:0] == 28'h000_0000, p3_reverse_8428_comb[27] && p3_reverse_8428_comb[26:0] == 27'h000_0000, p3_reverse_8428_comb[26] && p3_reverse_8428_comb[25:0] == 26'h000_0000, p3_reverse_8428_comb[25] && p3_reverse_8428_comb[24:0] == 25'h000_0000, p3_reverse_8428_comb[24] && p3_reverse_8428_comb[23:0] == 24'h00_0000, p3_reverse_8428_comb[23] && p3_reverse_8428_comb[22:0] == 23'h00_0000, p3_reverse_8428_comb[22] && p3_reverse_8428_comb[21:0] == 22'h00_0000, p3_reverse_8428_comb[21] && p3_reverse_8428_comb[20:0] == 21'h00_0000, p3_reverse_8428_comb[20] && p3_reverse_8428_comb[19:0] == 20'h0_0000, p3_reverse_8428_comb[19] && p3_reverse_8428_comb[18:0] == 19'h0_0000, p3_reverse_8428_comb[18] && p3_reverse_8428_comb[17:0] == 18'h0_0000, p3_reverse_8428_comb[17] && p3_reverse_8428_comb[16:0] == 17'h0_0000, p3_reverse_8428_comb[16] && p3_reverse_8428_comb[15:0] == 16'h0000, p3_reverse_8428_comb[15] && p3_reverse_8428_comb[14:0] == 15'h0000, p3_reverse_8428_comb[14] && p3_reverse_8428_comb[13:0] == 14'h0000, p3_reverse_8428_comb[13] && p3_reverse_8428_comb[12:0] == 13'h0000, p3_reverse_8428_comb[12] && p3_reverse_8428_comb[11:0] == 12'h000, p3_reverse_8428_comb[11] && p3_reverse_8428_comb[10:0] == 11'h000, p3_reverse_8428_comb[10] && p3_reverse_8428_comb[9:0] == 10'h000, p3_reverse_8428_comb[9] && p3_reverse_8428_comb[8:0] == 9'h000, p3_reverse_8428_comb[8] && p3_reverse_8428_comb[7:0] == 8'h00, p3_reverse_8428_comb[7] && p3_reverse_8428_comb[6:0] == 7'h00, p3_reverse_8428_comb[6] && p3_reverse_8428_comb[5:0] == 6'h00, p3_reverse_8428_comb[5] && p3_reverse_8428_comb[4:0] == 5'h00, p3_reverse_8428_comb[4] && p3_reverse_8428_comb[3:0] == 4'h0, p3_reverse_8428_comb[3] && p3_reverse_8428_comb[2:0] == 3'h0, p3_reverse_8428_comb[2] && p3_reverse_8428_comb[1:0] == 2'h0, p3_reverse_8428_comb[1] && !p3_reverse_8428_comb[0], p3_reverse_8428_comb[0]};
  assign p3_one_hot_8433_comb = {p3_reverse_8429_comb[27:0] == 28'h000_0000, p3_reverse_8429_comb[27] && p3_reverse_8429_comb[26:0] == 27'h000_0000, p3_reverse_8429_comb[26] && p3_reverse_8429_comb[25:0] == 26'h000_0000, p3_reverse_8429_comb[25] && p3_reverse_8429_comb[24:0] == 25'h000_0000, p3_reverse_8429_comb[24] && p3_reverse_8429_comb[23:0] == 24'h00_0000, p3_reverse_8429_comb[23] && p3_reverse_8429_comb[22:0] == 23'h00_0000, p3_reverse_8429_comb[22] && p3_reverse_8429_comb[21:0] == 22'h00_0000, p3_reverse_8429_comb[21] && p3_reverse_8429_comb[20:0] == 21'h00_0000, p3_reverse_8429_comb[20] && p3_reverse_8429_comb[19:0] == 20'h0_0000, p3_reverse_8429_comb[19] && p3_reverse_8429_comb[18:0] == 19'h0_0000, p3_reverse_8429_comb[18] && p3_reverse_8429_comb[17:0] == 18'h0_0000, p3_reverse_8429_comb[17] && p3_reverse_8429_comb[16:0] == 17'h0_0000, p3_reverse_8429_comb[16] && p3_reverse_8429_comb[15:0] == 16'h0000, p3_reverse_8429_comb[15] && p3_reverse_8429_comb[14:0] == 15'h0000, p3_reverse_8429_comb[14] && p3_reverse_8429_comb[13:0] == 14'h0000, p3_reverse_8429_comb[13] && p3_reverse_8429_comb[12:0] == 13'h0000, p3_reverse_8429_comb[12] && p3_reverse_8429_comb[11:0] == 12'h000, p3_reverse_8429_comb[11] && p3_reverse_8429_comb[10:0] == 11'h000, p3_reverse_8429_comb[10] && p3_reverse_8429_comb[9:0] == 10'h000, p3_reverse_8429_comb[9] && p3_reverse_8429_comb[8:0] == 9'h000, p3_reverse_8429_comb[8] && p3_reverse_8429_comb[7:0] == 8'h00, p3_reverse_8429_comb[7] && p3_reverse_8429_comb[6:0] == 7'h00, p3_reverse_8429_comb[6] && p3_reverse_8429_comb[5:0] == 6'h00, p3_reverse_8429_comb[5] && p3_reverse_8429_comb[4:0] == 5'h00, p3_reverse_8429_comb[4] && p3_reverse_8429_comb[3:0] == 4'h0, p3_reverse_8429_comb[3] && p3_reverse_8429_comb[2:0] == 3'h0, p3_reverse_8429_comb[2] && p3_reverse_8429_comb[1:0] == 2'h0, p3_reverse_8429_comb[1] && !p3_reverse_8429_comb[0], p3_reverse_8429_comb[0]};
  assign p3_one_hot_8434_comb = {p3_reverse_8430_comb[27:0] == 28'h000_0000, p3_reverse_8430_comb[27] && p3_reverse_8430_comb[26:0] == 27'h000_0000, p3_reverse_8430_comb[26] && p3_reverse_8430_comb[25:0] == 26'h000_0000, p3_reverse_8430_comb[25] && p3_reverse_8430_comb[24:0] == 25'h000_0000, p3_reverse_8430_comb[24] && p3_reverse_8430_comb[23:0] == 24'h00_0000, p3_reverse_8430_comb[23] && p3_reverse_8430_comb[22:0] == 23'h00_0000, p3_reverse_8430_comb[22] && p3_reverse_8430_comb[21:0] == 22'h00_0000, p3_reverse_8430_comb[21] && p3_reverse_8430_comb[20:0] == 21'h00_0000, p3_reverse_8430_comb[20] && p3_reverse_8430_comb[19:0] == 20'h0_0000, p3_reverse_8430_comb[19] && p3_reverse_8430_comb[18:0] == 19'h0_0000, p3_reverse_8430_comb[18] && p3_reverse_8430_comb[17:0] == 18'h0_0000, p3_reverse_8430_comb[17] && p3_reverse_8430_comb[16:0] == 17'h0_0000, p3_reverse_8430_comb[16] && p3_reverse_8430_comb[15:0] == 16'h0000, p3_reverse_8430_comb[15] && p3_reverse_8430_comb[14:0] == 15'h0000, p3_reverse_8430_comb[14] && p3_reverse_8430_comb[13:0] == 14'h0000, p3_reverse_8430_comb[13] && p3_reverse_8430_comb[12:0] == 13'h0000, p3_reverse_8430_comb[12] && p3_reverse_8430_comb[11:0] == 12'h000, p3_reverse_8430_comb[11] && p3_reverse_8430_comb[10:0] == 11'h000, p3_reverse_8430_comb[10] && p3_reverse_8430_comb[9:0] == 10'h000, p3_reverse_8430_comb[9] && p3_reverse_8430_comb[8:0] == 9'h000, p3_reverse_8430_comb[8] && p3_reverse_8430_comb[7:0] == 8'h00, p3_reverse_8430_comb[7] && p3_reverse_8430_comb[6:0] == 7'h00, p3_reverse_8430_comb[6] && p3_reverse_8430_comb[5:0] == 6'h00, p3_reverse_8430_comb[5] && p3_reverse_8430_comb[4:0] == 5'h00, p3_reverse_8430_comb[4] && p3_reverse_8430_comb[3:0] == 4'h0, p3_reverse_8430_comb[3] && p3_reverse_8430_comb[2:0] == 3'h0, p3_reverse_8430_comb[2] && p3_reverse_8430_comb[1:0] == 2'h0, p3_reverse_8430_comb[1] && !p3_reverse_8430_comb[0], p3_reverse_8430_comb[0]};
  assign p3_one_hot_8435_comb = {p3_reverse_8431_comb[27:0] == 28'h000_0000, p3_reverse_8431_comb[27] && p3_reverse_8431_comb[26:0] == 27'h000_0000, p3_reverse_8431_comb[26] && p3_reverse_8431_comb[25:0] == 26'h000_0000, p3_reverse_8431_comb[25] && p3_reverse_8431_comb[24:0] == 25'h000_0000, p3_reverse_8431_comb[24] && p3_reverse_8431_comb[23:0] == 24'h00_0000, p3_reverse_8431_comb[23] && p3_reverse_8431_comb[22:0] == 23'h00_0000, p3_reverse_8431_comb[22] && p3_reverse_8431_comb[21:0] == 22'h00_0000, p3_reverse_8431_comb[21] && p3_reverse_8431_comb[20:0] == 21'h00_0000, p3_reverse_8431_comb[20] && p3_reverse_8431_comb[19:0] == 20'h0_0000, p3_reverse_8431_comb[19] && p3_reverse_8431_comb[18:0] == 19'h0_0000, p3_reverse_8431_comb[18] && p3_reverse_8431_comb[17:0] == 18'h0_0000, p3_reverse_8431_comb[17] && p3_reverse_8431_comb[16:0] == 17'h0_0000, p3_reverse_8431_comb[16] && p3_reverse_8431_comb[15:0] == 16'h0000, p3_reverse_8431_comb[15] && p3_reverse_8431_comb[14:0] == 15'h0000, p3_reverse_8431_comb[14] && p3_reverse_8431_comb[13:0] == 14'h0000, p3_reverse_8431_comb[13] && p3_reverse_8431_comb[12:0] == 13'h0000, p3_reverse_8431_comb[12] && p3_reverse_8431_comb[11:0] == 12'h000, p3_reverse_8431_comb[11] && p3_reverse_8431_comb[10:0] == 11'h000, p3_reverse_8431_comb[10] && p3_reverse_8431_comb[9:0] == 10'h000, p3_reverse_8431_comb[9] && p3_reverse_8431_comb[8:0] == 9'h000, p3_reverse_8431_comb[8] && p3_reverse_8431_comb[7:0] == 8'h00, p3_reverse_8431_comb[7] && p3_reverse_8431_comb[6:0] == 7'h00, p3_reverse_8431_comb[6] && p3_reverse_8431_comb[5:0] == 6'h00, p3_reverse_8431_comb[5] && p3_reverse_8431_comb[4:0] == 5'h00, p3_reverse_8431_comb[4] && p3_reverse_8431_comb[3:0] == 4'h0, p3_reverse_8431_comb[3] && p3_reverse_8431_comb[2:0] == 3'h0, p3_reverse_8431_comb[2] && p3_reverse_8431_comb[1:0] == 2'h0, p3_reverse_8431_comb[1] && !p3_reverse_8431_comb[0], p3_reverse_8431_comb[0]};
  assign p3_encode_8436_comb = {p3_one_hot_8432_comb[16] | p3_one_hot_8432_comb[17] | p3_one_hot_8432_comb[18] | p3_one_hot_8432_comb[19] | p3_one_hot_8432_comb[20] | p3_one_hot_8432_comb[21] | p3_one_hot_8432_comb[22] | p3_one_hot_8432_comb[23] | p3_one_hot_8432_comb[24] | p3_one_hot_8432_comb[25] | p3_one_hot_8432_comb[26] | p3_one_hot_8432_comb[27] | p3_one_hot_8432_comb[28], p3_one_hot_8432_comb[8] | p3_one_hot_8432_comb[9] | p3_one_hot_8432_comb[10] | p3_one_hot_8432_comb[11] | p3_one_hot_8432_comb[12] | p3_one_hot_8432_comb[13] | p3_one_hot_8432_comb[14] | p3_one_hot_8432_comb[15] | p3_one_hot_8432_comb[24] | p3_one_hot_8432_comb[25] | p3_one_hot_8432_comb[26] | p3_one_hot_8432_comb[27] | p3_one_hot_8432_comb[28], p3_one_hot_8432_comb[4] | p3_one_hot_8432_comb[5] | p3_one_hot_8432_comb[6] | p3_one_hot_8432_comb[7] | p3_one_hot_8432_comb[12] | p3_one_hot_8432_comb[13] | p3_one_hot_8432_comb[14] | p3_one_hot_8432_comb[15] | p3_one_hot_8432_comb[20] | p3_one_hot_8432_comb[21] | p3_one_hot_8432_comb[22] | p3_one_hot_8432_comb[23] | p3_one_hot_8432_comb[28], p3_one_hot_8432_comb[2] | p3_one_hot_8432_comb[3] | p3_one_hot_8432_comb[6] | p3_one_hot_8432_comb[7] | p3_one_hot_8432_comb[10] | p3_one_hot_8432_comb[11] | p3_one_hot_8432_comb[14] | p3_one_hot_8432_comb[15] | p3_one_hot_8432_comb[18] | p3_one_hot_8432_comb[19] | p3_one_hot_8432_comb[22] | p3_one_hot_8432_comb[23] | p3_one_hot_8432_comb[26] | p3_one_hot_8432_comb[27], p3_one_hot_8432_comb[1] | p3_one_hot_8432_comb[3] | p3_one_hot_8432_comb[5] | p3_one_hot_8432_comb[7] | p3_one_hot_8432_comb[9] | p3_one_hot_8432_comb[11] | p3_one_hot_8432_comb[13] | p3_one_hot_8432_comb[15] | p3_one_hot_8432_comb[17] | p3_one_hot_8432_comb[19] | p3_one_hot_8432_comb[21] | p3_one_hot_8432_comb[23] | p3_one_hot_8432_comb[25] | p3_one_hot_8432_comb[27]};
  assign p3_encode_8437_comb = {p3_one_hot_8433_comb[16] | p3_one_hot_8433_comb[17] | p3_one_hot_8433_comb[18] | p3_one_hot_8433_comb[19] | p3_one_hot_8433_comb[20] | p3_one_hot_8433_comb[21] | p3_one_hot_8433_comb[22] | p3_one_hot_8433_comb[23] | p3_one_hot_8433_comb[24] | p3_one_hot_8433_comb[25] | p3_one_hot_8433_comb[26] | p3_one_hot_8433_comb[27] | p3_one_hot_8433_comb[28], p3_one_hot_8433_comb[8] | p3_one_hot_8433_comb[9] | p3_one_hot_8433_comb[10] | p3_one_hot_8433_comb[11] | p3_one_hot_8433_comb[12] | p3_one_hot_8433_comb[13] | p3_one_hot_8433_comb[14] | p3_one_hot_8433_comb[15] | p3_one_hot_8433_comb[24] | p3_one_hot_8433_comb[25] | p3_one_hot_8433_comb[26] | p3_one_hot_8433_comb[27] | p3_one_hot_8433_comb[28], p3_one_hot_8433_comb[4] | p3_one_hot_8433_comb[5] | p3_one_hot_8433_comb[6] | p3_one_hot_8433_comb[7] | p3_one_hot_8433_comb[12] | p3_one_hot_8433_comb[13] | p3_one_hot_8433_comb[14] | p3_one_hot_8433_comb[15] | p3_one_hot_8433_comb[20] | p3_one_hot_8433_comb[21] | p3_one_hot_8433_comb[22] | p3_one_hot_8433_comb[23] | p3_one_hot_8433_comb[28], p3_one_hot_8433_comb[2] | p3_one_hot_8433_comb[3] | p3_one_hot_8433_comb[6] | p3_one_hot_8433_comb[7] | p3_one_hot_8433_comb[10] | p3_one_hot_8433_comb[11] | p3_one_hot_8433_comb[14] | p3_one_hot_8433_comb[15] | p3_one_hot_8433_comb[18] | p3_one_hot_8433_comb[19] | p3_one_hot_8433_comb[22] | p3_one_hot_8433_comb[23] | p3_one_hot_8433_comb[26] | p3_one_hot_8433_comb[27], p3_one_hot_8433_comb[1] | p3_one_hot_8433_comb[3] | p3_one_hot_8433_comb[5] | p3_one_hot_8433_comb[7] | p3_one_hot_8433_comb[9] | p3_one_hot_8433_comb[11] | p3_one_hot_8433_comb[13] | p3_one_hot_8433_comb[15] | p3_one_hot_8433_comb[17] | p3_one_hot_8433_comb[19] | p3_one_hot_8433_comb[21] | p3_one_hot_8433_comb[23] | p3_one_hot_8433_comb[25] | p3_one_hot_8433_comb[27]};
  assign p3_encode_8438_comb = {p3_one_hot_8434_comb[16] | p3_one_hot_8434_comb[17] | p3_one_hot_8434_comb[18] | p3_one_hot_8434_comb[19] | p3_one_hot_8434_comb[20] | p3_one_hot_8434_comb[21] | p3_one_hot_8434_comb[22] | p3_one_hot_8434_comb[23] | p3_one_hot_8434_comb[24] | p3_one_hot_8434_comb[25] | p3_one_hot_8434_comb[26] | p3_one_hot_8434_comb[27] | p3_one_hot_8434_comb[28], p3_one_hot_8434_comb[8] | p3_one_hot_8434_comb[9] | p3_one_hot_8434_comb[10] | p3_one_hot_8434_comb[11] | p3_one_hot_8434_comb[12] | p3_one_hot_8434_comb[13] | p3_one_hot_8434_comb[14] | p3_one_hot_8434_comb[15] | p3_one_hot_8434_comb[24] | p3_one_hot_8434_comb[25] | p3_one_hot_8434_comb[26] | p3_one_hot_8434_comb[27] | p3_one_hot_8434_comb[28], p3_one_hot_8434_comb[4] | p3_one_hot_8434_comb[5] | p3_one_hot_8434_comb[6] | p3_one_hot_8434_comb[7] | p3_one_hot_8434_comb[12] | p3_one_hot_8434_comb[13] | p3_one_hot_8434_comb[14] | p3_one_hot_8434_comb[15] | p3_one_hot_8434_comb[20] | p3_one_hot_8434_comb[21] | p3_one_hot_8434_comb[22] | p3_one_hot_8434_comb[23] | p3_one_hot_8434_comb[28], p3_one_hot_8434_comb[2] | p3_one_hot_8434_comb[3] | p3_one_hot_8434_comb[6] | p3_one_hot_8434_comb[7] | p3_one_hot_8434_comb[10] | p3_one_hot_8434_comb[11] | p3_one_hot_8434_comb[14] | p3_one_hot_8434_comb[15] | p3_one_hot_8434_comb[18] | p3_one_hot_8434_comb[19] | p3_one_hot_8434_comb[22] | p3_one_hot_8434_comb[23] | p3_one_hot_8434_comb[26] | p3_one_hot_8434_comb[27], p3_one_hot_8434_comb[1] | p3_one_hot_8434_comb[3] | p3_one_hot_8434_comb[5] | p3_one_hot_8434_comb[7] | p3_one_hot_8434_comb[9] | p3_one_hot_8434_comb[11] | p3_one_hot_8434_comb[13] | p3_one_hot_8434_comb[15] | p3_one_hot_8434_comb[17] | p3_one_hot_8434_comb[19] | p3_one_hot_8434_comb[21] | p3_one_hot_8434_comb[23] | p3_one_hot_8434_comb[25] | p3_one_hot_8434_comb[27]};
  assign p3_encode_8439_comb = {p3_one_hot_8435_comb[16] | p3_one_hot_8435_comb[17] | p3_one_hot_8435_comb[18] | p3_one_hot_8435_comb[19] | p3_one_hot_8435_comb[20] | p3_one_hot_8435_comb[21] | p3_one_hot_8435_comb[22] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[24] | p3_one_hot_8435_comb[25] | p3_one_hot_8435_comb[26] | p3_one_hot_8435_comb[27] | p3_one_hot_8435_comb[28], p3_one_hot_8435_comb[8] | p3_one_hot_8435_comb[9] | p3_one_hot_8435_comb[10] | p3_one_hot_8435_comb[11] | p3_one_hot_8435_comb[12] | p3_one_hot_8435_comb[13] | p3_one_hot_8435_comb[14] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[24] | p3_one_hot_8435_comb[25] | p3_one_hot_8435_comb[26] | p3_one_hot_8435_comb[27] | p3_one_hot_8435_comb[28], p3_one_hot_8435_comb[4] | p3_one_hot_8435_comb[5] | p3_one_hot_8435_comb[6] | p3_one_hot_8435_comb[7] | p3_one_hot_8435_comb[12] | p3_one_hot_8435_comb[13] | p3_one_hot_8435_comb[14] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[20] | p3_one_hot_8435_comb[21] | p3_one_hot_8435_comb[22] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[28], p3_one_hot_8435_comb[2] | p3_one_hot_8435_comb[3] | p3_one_hot_8435_comb[6] | p3_one_hot_8435_comb[7] | p3_one_hot_8435_comb[10] | p3_one_hot_8435_comb[11] | p3_one_hot_8435_comb[14] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[18] | p3_one_hot_8435_comb[19] | p3_one_hot_8435_comb[22] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[26] | p3_one_hot_8435_comb[27], p3_one_hot_8435_comb[1] | p3_one_hot_8435_comb[3] | p3_one_hot_8435_comb[5] | p3_one_hot_8435_comb[7] | p3_one_hot_8435_comb[9] | p3_one_hot_8435_comb[11] | p3_one_hot_8435_comb[13] | p3_one_hot_8435_comb[15] | p3_one_hot_8435_comb[17] | p3_one_hot_8435_comb[19] | p3_one_hot_8435_comb[21] | p3_one_hot_8435_comb[23] | p3_one_hot_8435_comb[25] | p3_one_hot_8435_comb[27]};
  assign p3_carry_bit__2_comb = p3_abs_fraction__2_comb[27];
  assign p3_cancel__2_comb = p3_encode_8436_comb[1] | p3_encode_8436_comb[2] | p3_encode_8436_comb[3] | p3_encode_8436_comb[4];
  assign p3_carry_bit__3_comb = p3_abs_fraction__3_comb[27];
  assign p3_cancel__3_comb = p3_encode_8437_comb[1] | p3_encode_8437_comb[2] | p3_encode_8437_comb[3] | p3_encode_8437_comb[4];
  assign p3_carry_bit__4_comb = p3_abs_fraction__4_comb[27];
  assign p3_cancel__4_comb = p3_encode_8438_comb[1] | p3_encode_8438_comb[2] | p3_encode_8438_comb[3] | p3_encode_8438_comb[4];
  assign p3_carry_bit__5_comb = p3_abs_fraction__5_comb[27];
  assign p3_cancel__5_comb = p3_encode_8439_comb[1] | p3_encode_8439_comb[2] | p3_encode_8439_comb[3] | p3_encode_8439_comb[4];
  assign p3_leading_zeroes__2_comb = {23'h00_0000, p3_encode_8436_comb};
  assign p3_leading_zeroes__3_comb = {23'h00_0000, p3_encode_8437_comb};
  assign p3_leading_zeroes__4_comb = {23'h00_0000, p3_encode_8438_comb};
  assign p3_leading_zeroes__5_comb = {23'h00_0000, p3_encode_8439_comb};
  assign p3_carry_fraction__4_comb = p3_abs_fraction__2_comb[27:1];
  assign p3_add_8498_comb = p3_leading_zeroes__2_comb + 28'hfff_ffff;
  assign p3_carry_fraction__6_comb = p3_abs_fraction__3_comb[27:1];
  assign p3_add_8505_comb = p3_leading_zeroes__3_comb + 28'hfff_ffff;
  assign p3_carry_fraction__8_comb = p3_abs_fraction__4_comb[27:1];
  assign p3_add_8512_comb = p3_leading_zeroes__4_comb + 28'hfff_ffff;
  assign p3_carry_fraction__10_comb = p3_abs_fraction__5_comb[27:1];
  assign p3_add_8519_comb = p3_leading_zeroes__5_comb + 28'hfff_ffff;
  assign p3_concat_8520_comb = {~p3_carry_bit__2_comb & ~p3_cancel__2_comb, ~p3_carry_bit__2_comb & p3_cancel__2_comb, p3_carry_bit__2_comb & ~p3_cancel__2_comb};
  assign p3_carry_fraction__5_comb = p3_carry_fraction__4_comb | {26'h000_0000, p3_abs_fraction__2_comb[0]};
  assign p3_cancel_fraction__2_comb = p3_add_8498_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__2_comb[26:0] << p3_add_8498_comb;
  assign p3_concat_8523_comb = {~p3_carry_bit__3_comb & ~p3_cancel__3_comb, ~p3_carry_bit__3_comb & p3_cancel__3_comb, p3_carry_bit__3_comb & ~p3_cancel__3_comb};
  assign p3_carry_fraction__7_comb = p3_carry_fraction__6_comb | {26'h000_0000, p3_abs_fraction__3_comb[0]};
  assign p3_cancel_fraction__3_comb = p3_add_8505_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__3_comb[26:0] << p3_add_8505_comb;
  assign p3_concat_8526_comb = {~p3_carry_bit__4_comb & ~p3_cancel__4_comb, ~p3_carry_bit__4_comb & p3_cancel__4_comb, p3_carry_bit__4_comb & ~p3_cancel__4_comb};
  assign p3_carry_fraction__9_comb = p3_carry_fraction__8_comb | {26'h000_0000, p3_abs_fraction__4_comb[0]};
  assign p3_cancel_fraction__4_comb = p3_add_8512_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__4_comb[26:0] << p3_add_8512_comb;
  assign p3_concat_8529_comb = {~p3_carry_bit__5_comb & ~p3_cancel__5_comb, ~p3_carry_bit__5_comb & p3_cancel__5_comb, p3_carry_bit__5_comb & ~p3_cancel__5_comb};
  assign p3_carry_fraction__11_comb = p3_carry_fraction__10_comb | {26'h000_0000, p3_abs_fraction__5_comb[0]};
  assign p3_cancel_fraction__5_comb = p3_add_8519_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__5_comb[26:0] << p3_add_8519_comb;
  assign p3_shifted_fraction__2_comb = p3_carry_fraction__5_comb & {27{p3_concat_8520_comb[0]}} | p3_cancel_fraction__2_comb & {27{p3_concat_8520_comb[1]}} | p3_abs_fraction__2_comb[26:0] & {27{p3_concat_8520_comb[2]}};
  assign p3_shifted_fraction__3_comb = p3_carry_fraction__7_comb & {27{p3_concat_8523_comb[0]}} | p3_cancel_fraction__3_comb & {27{p3_concat_8523_comb[1]}} | p3_abs_fraction__3_comb[26:0] & {27{p3_concat_8523_comb[2]}};
  assign p3_shifted_fraction__4_comb = p3_carry_fraction__9_comb & {27{p3_concat_8526_comb[0]}} | p3_cancel_fraction__4_comb & {27{p3_concat_8526_comb[1]}} | p3_abs_fraction__4_comb[26:0] & {27{p3_concat_8526_comb[2]}};
  assign p3_shifted_fraction__5_comb = p3_carry_fraction__11_comb & {27{p3_concat_8529_comb[0]}} | p3_cancel_fraction__5_comb & {27{p3_concat_8529_comb[1]}} | p3_abs_fraction__5_comb[26:0] & {27{p3_concat_8529_comb[2]}};
  assign p3_normal_chunk__2_comb = p3_shifted_fraction__2_comb[2:0];
  assign p3_half_way_chunk__2_comb = p3_shifted_fraction__2_comb[3:2];
  assign p3_normal_chunk__3_comb = p3_shifted_fraction__3_comb[2:0];
  assign p3_half_way_chunk__3_comb = p3_shifted_fraction__3_comb[3:2];
  assign p3_normal_chunk__4_comb = p3_shifted_fraction__4_comb[2:0];
  assign p3_half_way_chunk__4_comb = p3_shifted_fraction__4_comb[3:2];
  assign p3_normal_chunk__5_comb = p3_shifted_fraction__5_comb[2:0];
  assign p3_half_way_chunk__5_comb = p3_shifted_fraction__5_comb[3:2];
  assign p3_add_8571_comb = {1'h0, p3_shifted_fraction__2_comb[26:3]} + 25'h000_0001;
  assign p3_add_8575_comb = {1'h0, p3_shifted_fraction__3_comb[26:3]} + 25'h000_0001;
  assign p3_add_8579_comb = {1'h0, p3_shifted_fraction__4_comb[26:3]} + 25'h000_0001;
  assign p3_add_8583_comb = {1'h0, p3_shifted_fraction__5_comb[26:3]} + 25'h000_0001;
  assign p3_do_round_up__7_comb = p3_normal_chunk__2_comb > 3'h4 | p3_half_way_chunk__2_comb == 2'h3;
  assign p3_do_round_up__8_comb = p3_normal_chunk__3_comb > 3'h4 | p3_half_way_chunk__3_comb == 2'h3;
  assign p3_do_round_up__9_comb = p3_normal_chunk__4_comb > 3'h4 | p3_half_way_chunk__4_comb == 2'h3;
  assign p3_do_round_up__10_comb = p3_normal_chunk__5_comb > 3'h4 | p3_half_way_chunk__5_comb == 2'h3;
  assign p3_rounded_fraction__2_comb = p3_do_round_up__7_comb ? {p3_add_8571_comb, p3_normal_chunk__2_comb} : {1'h0, p3_shifted_fraction__2_comb};
  assign p3_rounded_fraction__3_comb = p3_do_round_up__8_comb ? {p3_add_8575_comb, p3_normal_chunk__3_comb} : {1'h0, p3_shifted_fraction__3_comb};
  assign p3_rounded_fraction__4_comb = p3_do_round_up__9_comb ? {p3_add_8579_comb, p3_normal_chunk__4_comb} : {1'h0, p3_shifted_fraction__4_comb};
  assign p3_rounded_fraction__5_comb = p3_do_round_up__10_comb ? {p3_add_8583_comb, p3_normal_chunk__5_comb} : {1'h0, p3_shifted_fraction__5_comb};
  assign p3_rounding_carry__2_comb = p3_rounded_fraction__2_comb[27];
  assign p3_rounding_carry__3_comb = p3_rounded_fraction__3_comb[27];
  assign p3_rounding_carry__4_comb = p3_rounded_fraction__4_comb[27];
  assign p3_rounding_carry__5_comb = p3_rounded_fraction__5_comb[27];
  assign p3_concat_8610_comb = {1'h0, p2_greater_exp_bexp__2};
  assign p3_concat_8612_comb = {1'h0, p2_greater_exp_bexp__3};
  assign p3_add_8617_comb = p3_concat_8610_comb + {8'h00, p3_rounding_carry__2_comb};
  assign p3_add_8619_comb = p3_concat_8612_comb + {8'h00, p3_rounding_carry__3_comb};
  assign p3_add_8621_comb = p3_concat_8610_comb + {8'h00, p3_rounding_carry__4_comb};
  assign p3_add_8623_comb = p3_concat_8612_comb + {8'h00, p3_rounding_carry__5_comb};
  assign p3_add_8640_comb = {1'h0, p3_add_8617_comb} + 10'h001;
  assign p3_add_8643_comb = {1'h0, p3_add_8619_comb} + 10'h001;
  assign p3_add_8646_comb = {1'h0, p3_add_8621_comb} + 10'h001;
  assign p3_add_8649_comb = {1'h0, p3_add_8623_comb} + 10'h001;
  assign p3_wide_exponent__6_comb = p3_add_8640_comb - {5'h00, p3_encode_8436_comb};
  assign p3_wide_exponent__9_comb = p3_add_8643_comb - {5'h00, p3_encode_8437_comb};
  assign p3_wide_exponent__12_comb = p3_add_8646_comb - {5'h00, p3_encode_8438_comb};
  assign p3_wide_exponent__15_comb = p3_add_8649_comb - {5'h00, p3_encode_8439_comb};
  assign p3_wide_exponent__7_comb = p3_wide_exponent__6_comb & {10{p3_fraction__35_comb != 29'h0000_0000}};
  assign p3_wide_exponent__10_comb = p3_wide_exponent__9_comb & {10{p3_fraction__36_comb != 29'h0000_0000}};
  assign p3_wide_exponent__13_comb = p3_wide_exponent__12_comb & {10{p3_fraction__37_comb != 29'h0000_0000}};
  assign p3_wide_exponent__16_comb = p3_wide_exponent__15_comb & {10{p3_fraction__38_comb != 29'h0000_0000}};
  assign p3_wide_exponent__8_comb = p3_wide_exponent__7_comb[8:0] & {9{~p3_wide_exponent__7_comb[9]}};
  assign p3_wide_exponent__11_comb = p3_wide_exponent__10_comb[8:0] & {9{~p3_wide_exponent__10_comb[9]}};
  assign p3_wide_exponent__14_comb = p3_wide_exponent__13_comb[8:0] & {9{~p3_wide_exponent__13_comb[9]}};
  assign p3_wide_exponent__17_comb = p3_wide_exponent__16_comb[8:0] & {9{~p3_wide_exponent__16_comb[9]}};
  assign p3_fraction_is_zero__2_comb = p3_fraction__35_comb == 29'h0000_0000;
  assign p3_add_8744_comb = {2'h0, p3_rounding_carry__2_comb} + 3'h3;
  assign p3_fraction_is_zero__3_comb = p3_fraction__36_comb == 29'h0000_0000;
  assign p3_add_8750_comb = {2'h0, p3_rounding_carry__3_comb} + 3'h3;
  assign p3_fraction_is_zero__4_comb = p3_fraction__37_comb == 29'h0000_0000;
  assign p3_add_8756_comb = {2'h0, p3_rounding_carry__4_comb} + 3'h3;
  assign p3_fraction_is_zero__5_comb = p3_fraction__38_comb == 29'h0000_0000;
  assign p3_add_8762_comb = {2'h0, p3_rounding_carry__5_comb} + 3'h3;
  assign p3_nor_8766_comb = ~(p3_wide_exponent__8_comb[8] | p3_wide_exponent__8_comb[0] & p3_wide_exponent__8_comb[1] & p3_wide_exponent__8_comb[2] & p3_wide_exponent__8_comb[3] & p3_wide_exponent__8_comb[4] & p3_wide_exponent__8_comb[5] & p3_wide_exponent__8_comb[6] & p3_wide_exponent__8_comb[7]);
  assign p3_shrl_8767_comb = p3_rounded_fraction__2_comb >> p3_add_8744_comb;
  assign p3_nor_8771_comb = ~(p3_wide_exponent__11_comb[8] | p3_wide_exponent__11_comb[0] & p3_wide_exponent__11_comb[1] & p3_wide_exponent__11_comb[2] & p3_wide_exponent__11_comb[3] & p3_wide_exponent__11_comb[4] & p3_wide_exponent__11_comb[5] & p3_wide_exponent__11_comb[6] & p3_wide_exponent__11_comb[7]);
  assign p3_shrl_8772_comb = p3_rounded_fraction__3_comb >> p3_add_8750_comb;
  assign p3_nor_8776_comb = ~(p3_wide_exponent__14_comb[8] | p3_wide_exponent__14_comb[0] & p3_wide_exponent__14_comb[1] & p3_wide_exponent__14_comb[2] & p3_wide_exponent__14_comb[3] & p3_wide_exponent__14_comb[4] & p3_wide_exponent__14_comb[5] & p3_wide_exponent__14_comb[6] & p3_wide_exponent__14_comb[7]);
  assign p3_shrl_8777_comb = p3_rounded_fraction__4_comb >> p3_add_8756_comb;
  assign p3_nor_8781_comb = ~(p3_wide_exponent__17_comb[8] | p3_wide_exponent__17_comb[0] & p3_wide_exponent__17_comb[1] & p3_wide_exponent__17_comb[2] & p3_wide_exponent__17_comb[3] & p3_wide_exponent__17_comb[4] & p3_wide_exponent__17_comb[5] & p3_wide_exponent__17_comb[6] & p3_wide_exponent__17_comb[7]);
  assign p3_shrl_8782_comb = p3_rounded_fraction__5_comb >> p3_add_8762_comb;
  assign p3_result_sign__15_comb = ~(~p3_fraction__35_comb[28] | p3_greater_exp_sign__2_comb) | ~(p3_fraction__35_comb[28] | p3_fraction_is_zero__2_comb | ~p3_greater_exp_sign__2_comb);
  assign p3_result_fraction__19_comb = p3_shrl_8767_comb[22:0];
  assign p3_sign_ext_8789_comb = {23{p2_nor_8301}};
  assign p3_result_sign__17_comb = ~(~p3_fraction__36_comb[28] | p3_greater_exp_sign__3_comb) | ~(p3_fraction__36_comb[28] | p3_fraction_is_zero__3_comb | ~p3_greater_exp_sign__3_comb);
  assign p3_result_fraction__21_comb = p3_shrl_8772_comb[22:0];
  assign p3_sign_ext_8795_comb = {23{p2_nor_8305}};
  assign p3_result_sign__20_comb = ~(~p3_fraction__37_comb[28] | p3_greater_exp_sign__4_comb) | ~(p3_fraction__37_comb[28] | p3_fraction_is_zero__4_comb | ~p3_greater_exp_sign__4_comb);
  assign p3_result_fraction__24_comb = p3_shrl_8777_comb[22:0];
  assign p3_result_sign__23_comb = ~(~p3_fraction__38_comb[28] | p3_greater_exp_sign__5_comb) | ~(p3_fraction__38_comb[28] | p3_fraction_is_zero__5_comb | ~p3_greater_exp_sign__5_comb);
  assign p3_result_fraction__27_comb = p3_shrl_8782_comb[22:0];
  assign p3_result_sign__16_comb = p2_is_operand_inf__2 ? p2_not_8310 : p3_result_sign__15_comb;
  assign p3_high_exp__42_comb = 8'hff;
  assign p3_result_fraction__20_comb = p3_result_fraction__19_comb & {23{~(~(p3_wide_exponent__8_comb[1] | p3_wide_exponent__8_comb[2] | p3_wide_exponent__8_comb[3] | p3_wide_exponent__8_comb[4] | p3_wide_exponent__8_comb[5] | p3_wide_exponent__8_comb[6] | p3_wide_exponent__8_comb[7] | p3_wide_exponent__8_comb[8] | p3_wide_exponent__8_comb[0]))}} & {23{p3_nor_8766_comb}} & p3_sign_ext_8789_comb;
  assign p3_nan_fraction__16_comb = 23'h40_0000;
  assign p3_result_sign__18_comb = p2_is_operand_inf__3 ? p2_not_8313 : p3_result_sign__17_comb;
  assign p3_high_exp__43_comb = 8'hff;
  assign p3_result_fraction__22_comb = p3_result_fraction__21_comb & {23{~(~(p3_wide_exponent__11_comb[1] | p3_wide_exponent__11_comb[2] | p3_wide_exponent__11_comb[3] | p3_wide_exponent__11_comb[4] | p3_wide_exponent__11_comb[5] | p3_wide_exponent__11_comb[6] | p3_wide_exponent__11_comb[7] | p3_wide_exponent__11_comb[8] | p3_wide_exponent__11_comb[0]))}} & {23{p3_nor_8771_comb}} & p3_sign_ext_8795_comb;
  assign p3_nan_fraction__17_comb = 23'h40_0000;
  assign p3_result_sign__21_comb = p2_is_operand_inf__2 ? p2_not_8315 : p3_result_sign__20_comb;
  assign p3_high_exp__44_comb = 8'hff;
  assign p3_result_fraction__25_comb = p3_result_fraction__24_comb & {23{~(~(p3_wide_exponent__14_comb[1] | p3_wide_exponent__14_comb[2] | p3_wide_exponent__14_comb[3] | p3_wide_exponent__14_comb[4] | p3_wide_exponent__14_comb[5] | p3_wide_exponent__14_comb[6] | p3_wide_exponent__14_comb[7] | p3_wide_exponent__14_comb[8] | p3_wide_exponent__14_comb[0]))}} & {23{p3_nor_8776_comb}} & p3_sign_ext_8789_comb;
  assign p3_nan_fraction__18_comb = 23'h40_0000;
  assign p3_result_sign__24_comb = p2_is_operand_inf__3 ? p2_not_8317 : p3_result_sign__23_comb;
  assign p3_high_exp__45_comb = 8'hff;
  assign p3_result_fraction__28_comb = p3_result_fraction__27_comb & {23{~(~(p3_wide_exponent__17_comb[1] | p3_wide_exponent__17_comb[2] | p3_wide_exponent__17_comb[3] | p3_wide_exponent__17_comb[4] | p3_wide_exponent__17_comb[5] | p3_wide_exponent__17_comb[6] | p3_wide_exponent__17_comb[7] | p3_wide_exponent__17_comb[8] | p3_wide_exponent__17_comb[0]))}} & {23{p3_nor_8781_comb}} & p3_sign_ext_8795_comb;
  assign p3_nan_fraction__19_comb = 23'h40_0000;
  assign p3_result_sign__19_comb = ~p2_is_result_nan__7 & p3_result_sign__16_comb;
  assign p3_result_exponent__3_comb = p2_is_result_nan__7 | p2_is_operand_inf__2 | ~p3_nor_8766_comb ? p3_high_exp__42_comb : p3_wide_exponent__8_comb[7:0];
  assign p3_result_fraction__23_comb = p2_is_result_nan__7 ? p3_nan_fraction__16_comb : p3_result_fraction__20_comb;
  assign p3_result_sign__22_comb = ~p2_is_result_nan__8 & p3_result_sign__18_comb;
  assign p3_result_exponent__4_comb = p2_is_result_nan__8 | p2_is_operand_inf__3 | ~p3_nor_8771_comb ? p3_high_exp__43_comb : p3_wide_exponent__11_comb[7:0];
  assign p3_result_fraction__26_comb = p2_is_result_nan__8 ? p3_nan_fraction__17_comb : p3_result_fraction__22_comb;
  assign p3_result_sign__25_comb = ~p2_is_result_nan__9 & p3_result_sign__21_comb;
  assign p3_result_exponent__5_comb = p2_is_result_nan__9 | p2_is_operand_inf__2 | ~p3_nor_8776_comb ? p3_high_exp__44_comb : p3_wide_exponent__14_comb[7:0];
  assign p3_result_fraction__29_comb = p2_is_result_nan__9 ? p3_nan_fraction__18_comb : p3_result_fraction__25_comb;
  assign p3_result_sign__26_comb = ~p2_is_result_nan__10 & p3_result_sign__24_comb;
  assign p3_result_exponent__6_comb = p2_is_result_nan__10 | p2_is_operand_inf__3 | ~p3_nor_8781_comb ? p3_high_exp__45_comb : p3_wide_exponent__17_comb[7:0];
  assign p3_result_fraction__30_comb = p2_is_result_nan__10 ? p3_nan_fraction__19_comb : p3_result_fraction__28_comb;
  assign p3_out0_r_comb = {p3_result_sign__19_comb, p3_result_exponent__3_comb, p3_result_fraction__23_comb};
  assign p3_out0_i_comb = {p3_result_sign__22_comb, p3_result_exponent__4_comb, p3_result_fraction__26_comb};
  assign p3_out1_r_comb = {p3_result_sign__25_comb, p3_result_exponent__5_comb, p3_result_fraction__29_comb};
  assign p3_out1_i_comb = {p3_result_sign__26_comb, p3_result_exponent__6_comb, p3_result_fraction__30_comb};
  assign p3_tuple_8850_comb = {p3_out0_r_comb, p3_out0_i_comb, p3_out1_r_comb, p3_out1_i_comb};

  // Registers for pipe stage 3:
  reg [127:0] p3_tuple_8850;
  always_ff @ (posedge clk) begin
    p3_tuple_8850 <= p3_tuple_8850_comb;
  end
  assign out = p3_tuple_8850;
endmodule

module Neg #(
  parameter WIDTH = 32
) (
  input wire logic signed [WIDTH-1:0] in,
  output wire logic signed [WIDTH-1:0] out
);
  assign out = -in;
endmodule
`default_nettype none

module Register #(
    parameter WIDTH = 32
) (
  input wire clk,
  input wire reset,
  input wire logic write_en,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] out
);
  always_ff @(posedge clk) begin
    if (reset)
      out <= 0;
    else if (write_en)
      out <= in;
    else
      out <= out;
  end
endmodule

// Same as a register but does not have a write enable signal.
module Delay #(
    parameter WIDTH = 32
) (
  input wire clk,
  input wire reset,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] out
);

  Register #(WIDTH) r (
    .clk(clk),
    .reset(reset),
    .write_en(1'b1),
    .in(in),
    .out(out)
  );
endmodule

// Register that passes its input value through.
module PassThroughRegister #(
  parameter WIDTH = 32
) (
  input wire clk,
  input wire reset,
  input wire logic write_en,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] out
);
  // held register value
  logic [WIDTH-1:0] t_out;
  Register #(WIDTH) r (
    .clk(clk),
    .reset(reset),
    .write_en(write_en),
    .in(in),
    .out(t_out)
  );
  
  assign out = write_en ? in : t_out;
endmodule

// Similar to a register but provides access to its previous value only.
// Resetting behavior controlled using the SAFE parameter.
module Prev #(
    parameter WIDTH = 32,
    // If 0, reset to 'x, otherwise reset to 0
    parameter SAFE = 0
) (
  input wire clk,
  input wire reset,
  input wire logic write_en,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] prev
);
  always_ff @(posedge clk) begin
    if (reset)
      if (SAFE == 0)
        prev <= 'x;
      else
        prev <= '0;
    else if (write_en)
      prev <= in;
    else
      prev <= prev;
  end
endmodule

module ContPrev #(
    parameter WIDTH = 32,
    parameter SAFE = 0
) (
  input wire clk,
  input wire reset,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] prev
);

Prev #(WIDTH, SAFE) r (
  .clk(clk),
  .reset(reset),
  .write_en(1'b1),
  .in(in),
  .prev(prev)
);
endmodule


`default_nettype wire
module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module comp58(
  input logic [31:0] p2,
  output logic [31:0] p3,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp58
wire _guard0 = 1;
assign p3 = p2;
// COMPONENT END: comp58
endmodule
module comp60(
  input logic [31:0] p7,
  input logic [31:0] p8,
  output logic [63:0] p9,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp60
logic [31:0] inst0_p2;
logic [31:0] inst0_p3;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [31:0] inst1_right;
logic [63:0] inst1_out;
comp58 inst0 (
    .clk(inst0_clk),
    .p2(inst0_p2),
    .p3(inst0_p3),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(64),
    .RIGHT(32)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p9 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p3;
assign inst0_clk = clk;
assign inst0_p2 = p8;
assign inst0_reset = reset;
// COMPONENT END: comp60
endmodule
module comp61(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  output logic [95:0] p10,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp61
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [63:0] inst0_p9;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [63:0] inst1_right;
logic [95:0] inst1_out;
comp60 inst0 (
    .clk(inst0_clk),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(96),
    .RIGHT(64)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p10 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p9;
assign inst0_clk = clk;
assign inst0_p8 = p9;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp61
endmodule
module comp62(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  output logic [127:0] p11,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp62
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [95:0] inst0_p10;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [95:0] inst1_right;
logic [127:0] inst1_out;
comp61 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(128),
    .RIGHT(96)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p11 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p10;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p8 = p9;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp62
endmodule
module comp64(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  output logic [159:0] p12,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp64
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [127:0] inst0_p11;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [127:0] inst1_right;
logic [159:0] inst1_out;
comp62 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(160),
    .RIGHT(128)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p12 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p11;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp64
endmodule
module comp65(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  output logic [191:0] p13,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp65
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [159:0] inst0_p12;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [159:0] inst1_right;
logic [191:0] inst1_out;
comp64 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(192),
    .RIGHT(160)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p13 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p12;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp65
endmodule
module comp66(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  output logic [223:0] p14,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp66
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [191:0] inst0_p13;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [191:0] inst1_right;
logic [223:0] inst1_out;
comp65 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(224),
    .RIGHT(192)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p14 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p13;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp66
endmodule
module comp67(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  output logic [255:0] p15,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp67
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [223:0] inst0_p14;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [223:0] inst1_right;
logic [255:0] inst1_out;
comp66 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(256),
    .RIGHT(224)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p15 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p14;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
// COMPONENT END: comp67
endmodule
module comp68(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  output logic [287:0] p16,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp68
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [255:0] inst0_p15;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [255:0] inst1_right;
logic [287:0] inst1_out;
comp67 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(288),
    .RIGHT(256)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p16 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p15;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p14 = p15;
// COMPONENT END: comp68
endmodule
module comp69(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  output logic [319:0] p17,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp69
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [287:0] inst0_p16;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [287:0] inst1_right;
logic [319:0] inst1_out;
comp68 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(320),
    .RIGHT(288)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p17 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p16;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p14 = p15;
// COMPONENT END: comp69
endmodule
module comp70(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [351:0] p18,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp70
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [319:0] inst0_p17;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [319:0] inst1_right;
logic [351:0] inst1_out;
comp69 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(352),
    .RIGHT(320)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p18 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p17;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p14 = p15;
// COMPONENT END: comp70
endmodule
module comp71(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  output logic [383:0] p19,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp71
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [351:0] inst0_p18;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [351:0] inst1_right;
logic [383:0] inst1_out;
comp70 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(384),
    .RIGHT(352)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p19 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p18;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p14 = p15;
// COMPONENT END: comp71
endmodule
module comp72(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  output logic [415:0] p20,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp72
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [383:0] inst0_p19;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [383:0] inst1_right;
logic [415:0] inst1_out;
comp71 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(416),
    .RIGHT(384)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p20 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p19;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p14 = p15;
// COMPONENT END: comp72
endmodule
module comp73(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  output logic [447:0] p21,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp73
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [415:0] inst0_p20;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [415:0] inst1_right;
logic [447:0] inst1_out;
comp72 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(448),
    .RIGHT(416)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p21 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p20;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p14 = p15;
// COMPONENT END: comp73
endmodule
module comp74(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  output logic [479:0] p22,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp74
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [447:0] inst0_p21;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [447:0] inst1_right;
logic [479:0] inst1_out;
comp73 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(480),
    .RIGHT(448)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p22 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p21;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p14 = p15;
// COMPONENT END: comp74
endmodule
module comp75(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  output logic [511:0] p23,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp75
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [479:0] inst0_p22;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [479:0] inst1_right;
logic [511:0] inst1_out;
comp74 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(512),
    .RIGHT(480)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p23 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p22;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p14 = p15;
// COMPONENT END: comp75
endmodule
module comp76(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  output logic [543:0] p24,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp76
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [511:0] inst0_p23;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [511:0] inst1_right;
logic [543:0] inst1_out;
comp75 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(544),
    .RIGHT(512)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p24 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p23;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp76
endmodule
module comp77(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  output logic [575:0] p25,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp77
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [543:0] inst0_p24;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [543:0] inst1_right;
logic [575:0] inst1_out;
comp76 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(576),
    .RIGHT(544)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p25 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p24;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp77
endmodule
module comp78(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  output logic [607:0] p26,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp78
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [575:0] inst0_p25;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [575:0] inst1_right;
logic [607:0] inst1_out;
comp77 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(608),
    .RIGHT(576)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p26 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p25;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp78
endmodule
module comp79(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  output logic [639:0] p27,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp79
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [607:0] inst0_p26;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [607:0] inst1_right;
logic [639:0] inst1_out;
comp78 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(640),
    .RIGHT(608)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p27 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p26;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp79
endmodule
module comp80(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  output logic [671:0] p28,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp80
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [639:0] inst0_p27;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [639:0] inst1_right;
logic [671:0] inst1_out;
comp79 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(672),
    .RIGHT(640)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p28 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p27;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p22 = p23;
// COMPONENT END: comp80
endmodule
module comp81(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  output logic [703:0] p29,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp81
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [671:0] inst0_p28;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [671:0] inst1_right;
logic [703:0] inst1_out;
comp80 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(704),
    .RIGHT(672)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p29 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p28;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp81
endmodule
module comp53(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp53
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p10;
assign p29 = p11;
assign p20 = p2;
assign p21 = p3;
assign p23 = p3;
assign p25 = p3;
assign p18 = p2;
assign p30 = p10;
assign p24 = p2;
assign p32 = p10;
assign p26 = p10;
assign p31 = p11;
assign p27 = p11;
assign p33 = p11;
assign p22 = p2;
// COMPONENT END: comp53
endmodule
module comp42(
  output logic [31:0] p2,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp42
logic [31:0] inst0_out;
Const # (
    .VALUE(1060439283),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp42
endmodule
module comp39(
  output logic [31:0] p2,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp39
logic [31:0] inst0_out;
Const # (
    .VALUE(1064076126),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp39
endmodule
module comp82(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  output logic [735:0] p30,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp82
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [703:0] inst0_p29;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [703:0] inst1_right;
logic [735:0] inst1_out;
comp81 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(736),
    .RIGHT(704)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p30 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p29;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp82
endmodule
module comp83(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  output logic [767:0] p31,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp83
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [735:0] inst0_p30;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [735:0] inst1_right;
logic [767:0] inst1_out;
comp82 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(768),
    .RIGHT(736)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p31 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p30;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp83
endmodule
module comp84(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  output logic [799:0] p32,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp84
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [767:0] inst0_p31;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [767:0] inst1_right;
logic [799:0] inst1_out;
comp83 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(800),
    .RIGHT(768)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p32 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p31;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp84
endmodule
module comp85(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  output logic [831:0] p33,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp85
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [799:0] inst0_p32;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [799:0] inst1_right;
logic [831:0] inst1_out;
comp84 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(832),
    .RIGHT(800)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p33 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p32;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp85
endmodule
module comp86(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  output logic [863:0] p34,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp86
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [831:0] inst0_p33;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [831:0] inst1_right;
logic [863:0] inst1_out;
comp85 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(864),
    .RIGHT(832)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p34 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p33;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp86
endmodule
module comp87(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  output logic [895:0] p35,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp87
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [863:0] inst0_p34;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [863:0] inst1_right;
logic [895:0] inst1_out;
comp86 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(896),
    .RIGHT(864)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p35 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p34;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
// COMPONENT END: comp87
endmodule
module comp88(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  output logic [927:0] p36,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp88
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [895:0] inst0_p35;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [895:0] inst1_right;
logic [927:0] inst1_out;
comp87 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(928),
    .RIGHT(896)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p36 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p35;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
// COMPONENT END: comp88
endmodule
module comp89(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  output logic [959:0] p37,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp89
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [927:0] inst0_p36;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [927:0] inst1_right;
logic [959:0] inst1_out;
comp88 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(960),
    .RIGHT(928)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p37 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p36;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
assign inst0_p35 = p36;
// COMPONENT END: comp89
endmodule
module comp90(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  input logic [31:0] p37,
  output logic [991:0] p38,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp90
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [959:0] inst0_p37;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [959:0] inst1_right;
logic [991:0] inst1_out;
comp89 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(992),
    .RIGHT(960)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p38 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p37;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p36 = p37;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
assign inst0_p35 = p36;
// COMPONENT END: comp90
endmodule
module comp91(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  input logic [31:0] p37,
  input logic [31:0] p38,
  output logic [1023:0] p39,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp91
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [991:0] inst0_p38;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [991:0] inst1_right;
logic [1023:0] inst1_out;
comp90 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(1024),
    .RIGHT(992)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p39 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p38;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p36 = p37;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
assign inst0_p35 = p36;
assign inst0_p37 = p38;
// COMPONENT END: comp91
endmodule
module comp1(
  input logic [31:0] p2,
  output logic [31:0] p3,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp1
wire _guard0 = 1;
assign p3 = p2;
// COMPONENT END: comp1
endmodule
module comp2(
  input logic [63:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp2
logic [63:0] inst0_in;
logic [31:0] inst0_out;
logic [63:0] inst1_in;
logic [31:0] inst1_out;
logic [31:0] inst2_p2;
logic [31:0] inst2_p3;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(64),
    .LSB(32),
    .MSB(63),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(64),
    .LSB(0),
    .MSB(31),
    .OUT_WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp1 inst2 (
    .clk(inst2_clk),
    .p2(inst2_p2),
    .p3(inst2_p3),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p9 = inst0_out;
assign p10 = inst2_p3;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p2 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp2
endmodule
module comp3(
  input logic [95:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp3
logic [95:0] inst0_in;
logic [31:0] inst0_out;
logic [95:0] inst1_in;
logic [63:0] inst1_out;
logic [63:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(96),
    .LSB(64),
    .MSB(95),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(96),
    .LSB(0),
    .MSB(63),
    .OUT_WIDTH(64)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp2 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp3
endmodule
module comp4(
  input logic [127:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp4
logic [127:0] inst0_in;
logic [31:0] inst0_out;
logic [127:0] inst1_in;
logic [95:0] inst1_out;
logic [95:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(128),
    .LSB(96),
    .MSB(127),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(0),
    .MSB(95),
    .OUT_WIDTH(96)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp3 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp4
endmodule
module comp5(
  input logic [159:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp5
logic [159:0] inst0_in;
logic [31:0] inst0_out;
logic [159:0] inst1_in;
logic [127:0] inst1_out;
logic [127:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(160),
    .LSB(128),
    .MSB(159),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(160),
    .LSB(0),
    .MSB(127),
    .OUT_WIDTH(128)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp4 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp5
endmodule
module comp6(
  input logic [191:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp6
logic [191:0] inst0_in;
logic [31:0] inst0_out;
logic [191:0] inst1_in;
logic [159:0] inst1_out;
logic [159:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(192),
    .LSB(160),
    .MSB(191),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(192),
    .LSB(0),
    .MSB(159),
    .OUT_WIDTH(160)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp5 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp6
endmodule
module comp7(
  input logic [223:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp7
logic [223:0] inst0_in;
logic [31:0] inst0_out;
logic [223:0] inst1_in;
logic [191:0] inst1_out;
logic [191:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(224),
    .LSB(192),
    .MSB(223),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(224),
    .LSB(0),
    .MSB(191),
    .OUT_WIDTH(192)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp6 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp7
endmodule
module comp8(
  input logic [255:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp8
logic [255:0] inst0_in;
logic [31:0] inst0_out;
logic [255:0] inst1_in;
logic [223:0] inst1_out;
logic [223:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(256),
    .LSB(224),
    .MSB(255),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(256),
    .LSB(0),
    .MSB(223),
    .OUT_WIDTH(224)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp7 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp8
endmodule
module comp9(
  input logic [287:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp9
logic [287:0] inst0_in;
logic [31:0] inst0_out;
logic [287:0] inst1_in;
logic [255:0] inst1_out;
logic [255:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(288),
    .LSB(256),
    .MSB(287),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(288),
    .LSB(0),
    .MSB(255),
    .OUT_WIDTH(256)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp8 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp9
endmodule
module comp10(
  input logic [319:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp10
logic [319:0] inst0_in;
logic [31:0] inst0_out;
logic [319:0] inst1_in;
logic [287:0] inst1_out;
logic [287:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(320),
    .LSB(288),
    .MSB(319),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(320),
    .LSB(0),
    .MSB(287),
    .OUT_WIDTH(288)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp9 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp10
endmodule
module comp11(
  input logic [351:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp11
logic [351:0] inst0_in;
logic [31:0] inst0_out;
logic [351:0] inst1_in;
logic [319:0] inst1_out;
logic [319:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(352),
    .LSB(320),
    .MSB(351),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(352),
    .LSB(0),
    .MSB(319),
    .OUT_WIDTH(320)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp10 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp11
endmodule
module comp12(
  input logic [383:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp12
logic [383:0] inst0_in;
logic [31:0] inst0_out;
logic [383:0] inst1_in;
logic [351:0] inst1_out;
logic [351:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(384),
    .LSB(352),
    .MSB(383),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(384),
    .LSB(0),
    .MSB(351),
    .OUT_WIDTH(352)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp11 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp12
endmodule
module comp13(
  input logic [415:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp13
logic [415:0] inst0_in;
logic [31:0] inst0_out;
logic [415:0] inst1_in;
logic [383:0] inst1_out;
logic [383:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(416),
    .LSB(384),
    .MSB(415),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(416),
    .LSB(0),
    .MSB(383),
    .OUT_WIDTH(384)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp12 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp13
endmodule
module comp14(
  input logic [447:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp14
logic [447:0] inst0_in;
logic [31:0] inst0_out;
logic [447:0] inst1_in;
logic [415:0] inst1_out;
logic [415:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(448),
    .LSB(416),
    .MSB(447),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(448),
    .LSB(0),
    .MSB(415),
    .OUT_WIDTH(416)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp13 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp14
endmodule
module comp15(
  input logic [479:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp15
logic [479:0] inst0_in;
logic [31:0] inst0_out;
logic [479:0] inst1_in;
logic [447:0] inst1_out;
logic [447:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(480),
    .LSB(448),
    .MSB(479),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(480),
    .LSB(0),
    .MSB(447),
    .OUT_WIDTH(448)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp14 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp15
endmodule
module comp16(
  input logic [511:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp16
logic [511:0] inst0_in;
logic [31:0] inst0_out;
logic [511:0] inst1_in;
logic [479:0] inst1_out;
logic [479:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(512),
    .LSB(480),
    .MSB(511),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(512),
    .LSB(0),
    .MSB(479),
    .OUT_WIDTH(480)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp15 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp16
endmodule
module comp17(
  input logic [543:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp17
logic [543:0] inst0_in;
logic [31:0] inst0_out;
logic [543:0] inst1_in;
logic [511:0] inst1_out;
logic [511:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(544),
    .LSB(512),
    .MSB(543),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(544),
    .LSB(0),
    .MSB(511),
    .OUT_WIDTH(512)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp16 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp17
endmodule
module comp18(
  input logic [575:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp18
logic [575:0] inst0_in;
logic [31:0] inst0_out;
logic [575:0] inst1_in;
logic [543:0] inst1_out;
logic [543:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(576),
    .LSB(544),
    .MSB(575),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(576),
    .LSB(0),
    .MSB(543),
    .OUT_WIDTH(544)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp17 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp18
endmodule
module comp38(
  output logic [31:0] p2,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp38
logic [31:0] inst0_out;
Const # (
    .VALUE(621621554),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp38
endmodule
module comp46(
  output logic [31:0] p2,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp46
logic [31:0] inst0_out;
Const # (
    .VALUE(613232946),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp46
endmodule
module comp37(
  output logic [31:0] p2,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp37
logic [31:0] inst0_out;
Const # (
    .VALUE(1065353216),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp37
endmodule
module comp45(
  output logic [31:0] p4,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp45
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1083407522),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp45
endmodule
module comp47(
  output logic [31:0] p4,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp47
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1082130432),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp47
endmodule
module comp43(
  output logic [31:0] p4,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp43
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1087044365),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp43
endmodule
module comp41(
  output logic [31:0] p4,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp41
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1094455531),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp41
endmodule
module comp44(
  output logic [31:0] p2,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp44
logic [31:0] inst0_out;
Const # (
    .VALUE(1053028117),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp44
endmodule
module comp48(
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp48
logic [31:0] inst0_p2;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_p2;
logic inst1_reset;
logic inst1_clk;
logic [31:0] inst2_p2;
logic inst2_reset;
logic inst2_clk;
logic [31:0] inst3_p4;
logic inst3_clk;
logic inst3_reset;
logic [31:0] inst4_p2;
logic inst4_clk;
logic inst4_reset;
logic [31:0] inst5_p4;
logic inst5_clk;
logic inst5_reset;
logic [31:0] inst6_p2;
logic inst6_reset;
logic inst6_clk;
logic [31:0] inst7_p4;
logic inst7_clk;
logic inst7_reset;
logic [31:0] inst8_p2;
logic inst8_clk;
logic inst8_reset;
logic [31:0] inst9_p4;
logic inst9_reset;
logic inst9_clk;
logic [31:0] inst10_p4;
logic inst10_clk;
logic inst10_reset;
logic [31:0] inst11_p4;
logic inst11_clk;
logic inst11_reset;
logic [31:0] inst12_p4;
logic inst12_clk;
logic inst12_reset;
logic [31:0] inst13_p4;
logic inst13_clk;
logic inst13_reset;
logic [31:0] inst14_p4;
logic inst14_clk;
logic inst14_reset;
logic [31:0] inst15_p4;
logic inst15_clk;
logic inst15_reset;
comp37 inst0 (
    .clk(inst0_clk),
    .p2(inst0_p2),
    .reset(inst0_reset)
);
comp38 inst1 (
    .clk(inst1_clk),
    .p2(inst1_p2),
    .reset(inst1_reset)
);
comp39 inst2 (
    .clk(inst2_clk),
    .p2(inst2_p2),
    .reset(inst2_reset)
);
comp41 inst3 (
    .clk(inst3_clk),
    .p4(inst3_p4),
    .reset(inst3_reset)
);
comp42 inst4 (
    .clk(inst4_clk),
    .p2(inst4_p2),
    .reset(inst4_reset)
);
comp43 inst5 (
    .clk(inst5_clk),
    .p4(inst5_p4),
    .reset(inst5_reset)
);
comp44 inst6 (
    .clk(inst6_clk),
    .p2(inst6_p2),
    .reset(inst6_reset)
);
comp45 inst7 (
    .clk(inst7_clk),
    .p4(inst7_p4),
    .reset(inst7_reset)
);
comp46 inst8 (
    .clk(inst8_clk),
    .p2(inst8_p2),
    .reset(inst8_reset)
);
comp47 inst9 (
    .clk(inst9_clk),
    .p4(inst9_p4),
    .reset(inst9_reset)
);
comp41 inst10 (
    .clk(inst10_clk),
    .p4(inst10_p4),
    .reset(inst10_reset)
);
comp45 inst11 (
    .clk(inst11_clk),
    .p4(inst11_p4),
    .reset(inst11_reset)
);
comp43 inst12 (
    .clk(inst12_clk),
    .p4(inst12_p4),
    .reset(inst12_reset)
);
comp43 inst13 (
    .clk(inst13_clk),
    .p4(inst13_p4),
    .reset(inst13_reset)
);
comp45 inst14 (
    .clk(inst14_clk),
    .p4(inst14_p4),
    .reset(inst14_reset)
);
comp41 inst15 (
    .clk(inst15_clk),
    .p4(inst15_p4),
    .reset(inst15_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p2;
assign p28 = inst11_p4;
assign p29 = inst12_p4;
assign p17 = inst0_p2;
assign p20 = inst3_p4;
assign p21 = inst4_p2;
assign p23 = inst6_p2;
assign p25 = inst8_p2;
assign p18 = inst1_p2;
assign p30 = inst13_p4;
assign p24 = inst7_p4;
assign p32 = inst15_p4;
assign p26 = inst9_p4;
assign p31 = inst14_p4;
assign p27 = inst10_p4;
assign p22 = inst5_p4;
assign inst5_clk = clk;
assign inst5_reset = reset;
assign inst15_clk = clk;
assign inst15_reset = reset;
assign inst8_clk = clk;
assign inst8_reset = reset;
assign inst12_clk = clk;
assign inst12_reset = reset;
assign inst3_clk = clk;
assign inst3_reset = reset;
assign inst9_clk = clk;
assign inst9_reset = reset;
assign inst1_clk = clk;
assign inst1_reset = reset;
assign inst0_clk = clk;
assign inst0_reset = reset;
assign inst7_clk = clk;
assign inst7_reset = reset;
assign inst6_clk = clk;
assign inst6_reset = reset;
assign inst14_clk = clk;
assign inst14_reset = reset;
assign inst2_clk = clk;
assign inst2_reset = reset;
assign inst4_clk = clk;
assign inst4_reset = reset;
assign inst10_clk = clk;
assign inst10_reset = reset;
assign inst11_clk = clk;
assign inst11_reset = reset;
assign inst13_clk = clk;
assign inst13_reset = reset;
// COMPONENT END: comp48
endmodule
module comp19(
  input logic [607:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp19
logic [607:0] inst0_in;
logic [31:0] inst0_out;
logic [607:0] inst1_in;
logic [575:0] inst1_out;
logic [575:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(608),
    .LSB(576),
    .MSB(607),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(608),
    .LSB(0),
    .MSB(575),
    .OUT_WIDTH(576)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp18 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp19
endmodule
module comp20(
  input logic [639:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp20
logic [639:0] inst0_in;
logic [31:0] inst0_out;
logic [639:0] inst1_in;
logic [607:0] inst1_out;
logic [607:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(640),
    .LSB(608),
    .MSB(639),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(640),
    .LSB(0),
    .MSB(607),
    .OUT_WIDTH(608)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp19 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp20
endmodule
module comp21(
  input logic [671:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp21
logic [671:0] inst0_in;
logic [31:0] inst0_out;
logic [671:0] inst1_in;
logic [639:0] inst1_out;
logic [639:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(672),
    .LSB(640),
    .MSB(671),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(672),
    .LSB(0),
    .MSB(639),
    .OUT_WIDTH(640)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp20 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp21
endmodule
module comp22(
  input logic [703:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp22
logic [703:0] inst0_in;
logic [31:0] inst0_out;
logic [703:0] inst1_in;
logic [671:0] inst1_out;
logic [671:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(704),
    .LSB(672),
    .MSB(703),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(704),
    .LSB(0),
    .MSB(671),
    .OUT_WIDTH(672)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp21 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp22
endmodule
module comp23(
  input logic [735:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp23
logic [735:0] inst0_in;
logic [31:0] inst0_out;
logic [735:0] inst1_in;
logic [703:0] inst1_out;
logic [703:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(736),
    .LSB(704),
    .MSB(735),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(736),
    .LSB(0),
    .MSB(703),
    .OUT_WIDTH(704)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp22 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp23
endmodule
module comp24(
  input logic [767:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp24
logic [767:0] inst0_in;
logic [31:0] inst0_out;
logic [767:0] inst1_in;
logic [735:0] inst1_out;
logic [735:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(768),
    .LSB(736),
    .MSB(767),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(768),
    .LSB(0),
    .MSB(735),
    .OUT_WIDTH(736)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp23 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp24
endmodule
module comp25(
  input logic [799:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp25
logic [799:0] inst0_in;
logic [31:0] inst0_out;
logic [799:0] inst1_in;
logic [767:0] inst1_out;
logic [767:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(800),
    .LSB(768),
    .MSB(799),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(800),
    .LSB(0),
    .MSB(767),
    .OUT_WIDTH(768)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp24 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp25
endmodule
module comp26(
  input logic [831:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp26
logic [831:0] inst0_in;
logic [31:0] inst0_out;
logic [831:0] inst1_in;
logic [799:0] inst1_out;
logic [799:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(832),
    .LSB(800),
    .MSB(831),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(832),
    .LSB(0),
    .MSB(799),
    .OUT_WIDTH(800)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp25 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp26
endmodule
module comp27(
  input logic [863:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp27
logic [863:0] inst0_in;
logic [31:0] inst0_out;
logic [863:0] inst1_in;
logic [831:0] inst1_out;
logic [831:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(864),
    .LSB(832),
    .MSB(863),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(864),
    .LSB(0),
    .MSB(831),
    .OUT_WIDTH(832)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp26 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp27
endmodule
module comp28(
  input logic [895:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp28
logic [895:0] inst0_in;
logic [31:0] inst0_out;
logic [895:0] inst1_in;
logic [863:0] inst1_out;
logic [863:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(896),
    .LSB(864),
    .MSB(895),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(896),
    .LSB(0),
    .MSB(863),
    .OUT_WIDTH(864)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp27 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp28
endmodule
module comp29(
  input logic [927:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp29
logic [927:0] inst0_in;
logic [31:0] inst0_out;
logic [927:0] inst1_in;
logic [895:0] inst1_out;
logic [895:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(928),
    .LSB(896),
    .MSB(927),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(928),
    .LSB(0),
    .MSB(895),
    .OUT_WIDTH(896)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp28 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp29
endmodule
module comp30(
  input logic [959:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp30
logic [959:0] inst0_in;
logic [31:0] inst0_out;
logic [959:0] inst1_in;
logic [927:0] inst1_out;
logic [927:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(960),
    .LSB(928),
    .MSB(959),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(960),
    .LSB(0),
    .MSB(927),
    .OUT_WIDTH(928)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp29 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p38 = inst2_p37;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp30
endmodule
module comp50(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  output logic [31:0] p40,
  output logic [31:0] p41,
  output logic [31:0] p42,
  output logic [31:0] p43,
  output logic [31:0] p44,
  output logic [31:0] p45,
  output logic [31:0] p46,
  output logic [31:0] p47,
  output logic [31:0] p48,
  output logic [31:0] p49,
  output logic [31:0] p50,
  output logic [31:0] p51,
  output logic [31:0] p52,
  output logic [31:0] p53,
  output logic [31:0] p54,
  output logic [31:0] p55,
  output logic [31:0] p56,
  output logic [31:0] p57,
  output logic [31:0] p58,
  output logic [31:0] p59,
  output logic [31:0] p60,
  output logic [31:0] p61,
  output logic [31:0] p62,
  output logic [31:0] p63,
  output logic [31:0] p64,
  output logic [31:0] p65,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp50
wire _guard0 = 1;
assign p38 = p10;
assign p40 = p26;
assign p47 = p15;
assign p65 = p33;
assign p52 = p20;
assign p59 = p9;
assign p56 = p28;
assign p60 = p24;
assign p64 = p32;
assign p36 = p18;
assign p39 = p11;
assign p46 = p14;
assign p51 = p5;
assign p54 = p12;
assign p45 = p23;
assign p53 = p21;
assign p58 = p8;
assign p50 = p4;
assign p41 = p27;
assign p43 = p7;
assign p63 = p17;
assign p42 = p6;
assign p48 = p30;
assign p49 = p31;
assign p61 = p25;
assign p62 = p16;
assign p34 = p2;
assign p35 = p3;
assign p57 = p29;
assign p37 = p19;
assign p44 = p22;
assign p55 = p13;
// COMPONENT END: comp50
endmodule
module comp52(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp52
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p2;
assign p29 = p3;
assign p20 = p2;
assign p21 = p3;
assign p23 = p3;
assign p25 = p3;
assign p18 = p2;
assign p30 = p2;
assign p24 = p2;
assign p32 = p2;
assign p26 = p2;
assign p31 = p3;
assign p27 = p3;
assign p33 = p3;
assign p22 = p2;
// COMPONENT END: comp52
endmodule
module comp34(
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp34
logic [31:0] inst0_in0_r;
logic [31:0] inst0_in0_i;
logic [31:0] inst0_in1_r;
logic [31:0] inst0_in1_i;
logic [31:0] inst0_twd_r;
logic [31:0] inst0_twd_i;
logic [127:0] inst0_out;
logic inst0_clk;
logic [127:0] inst1_in;
logic [31:0] inst1_out;
logic [127:0] inst2_in;
logic [31:0] inst2_out;
logic [127:0] inst3_in;
logic [31:0] inst3_out;
logic [127:0] inst4_in;
logic [31:0] inst4_out;
Butterfly_Exp8_Mant23 inst0 (
    .clk(inst0_clk),
    .in0_i(inst0_in0_i),
    .in0_r(inst0_in0_r),
    .in1_i(inst0_in1_i),
    .in1_r(inst0_in1_r),
    .out(inst0_out),
    .twd_i(inst0_twd_i),
    .twd_r(inst0_twd_r)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(96),
    .MSB(127),
    .OUT_WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(64),
    .MSB(95),
    .OUT_WIDTH(32)
) inst2 (
    .in(inst2_in),
    .out(inst2_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(32),
    .MSB(63),
    .OUT_WIDTH(32)
) inst3 (
    .in(inst3_in),
    .out(inst3_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(0),
    .MSB(31),
    .OUT_WIDTH(32)
) inst4 (
    .in(inst4_in),
    .out(inst4_out)
);
wire _guard0 = 1;
assign p28 = inst3_out;
assign p29 = inst4_out;
assign p26 = inst1_out;
assign p27 = inst2_out;
assign inst3_in = inst0_out;
assign inst1_in = inst0_out;
assign inst0_in1_i = p23;
assign inst0_twd_i = p25;
assign inst0_clk = clk;
assign inst0_in0_i = p21;
assign inst0_in1_r = p22;
assign inst0_twd_r = p24;
assign inst0_in0_r = p20;
assign inst2_in = inst0_out;
assign inst4_in = inst0_out;
// COMPONENT END: comp34
endmodule
module comp31(
  input logic [991:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp31
logic [991:0] inst0_in;
logic [31:0] inst0_out;
logic [991:0] inst1_in;
logic [959:0] inst1_out;
logic [959:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic [31:0] inst2_p38;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(992),
    .LSB(960),
    .MSB(991),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(992),
    .LSB(0),
    .MSB(959),
    .OUT_WIDTH(960)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp30 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p38(inst2_p38),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p38 = inst2_p37;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p39 = inst2_p38;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp31
endmodule
module comp32(
  input logic [1023:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  output logic [31:0] p40,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp32
logic [1023:0] inst0_in;
logic [31:0] inst0_out;
logic [1023:0] inst1_in;
logic [991:0] inst1_out;
logic [991:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic [31:0] inst2_p38;
logic [31:0] inst2_p39;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(1024),
    .LSB(992),
    .MSB(1023),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(1024),
    .LSB(0),
    .MSB(991),
    .OUT_WIDTH(992)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp31 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p38(inst2_p38),
    .p39(inst2_p39),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p38 = inst2_p37;
assign p40 = inst2_p39;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p39 = inst2_p38;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp32
endmodule
module comp93(
  input logic [1023:0] p4,
  output logic [31:0] p5,
  output logic [31:0] p6,
  output logic [31:0] p7,
  output logic [31:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp93
logic [1023:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [31:0] inst0_p38;
logic [31:0] inst0_p39;
logic [31:0] inst0_p40;
logic inst0_reset;
logic inst0_clk;
comp32 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p39(inst0_p39),
    .p40(inst0_p40),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
wire _guard0 = 1;
assign p19 = inst0_p23;
assign p28 = inst0_p32;
assign p29 = inst0_p33;
assign p12 = inst0_p16;
assign p16 = inst0_p20;
assign p6 = inst0_p10;
assign p9 = inst0_p13;
assign p15 = inst0_p19;
assign p17 = inst0_p21;
assign p20 = inst0_p24;
assign p21 = inst0_p25;
assign p23 = inst0_p27;
assign p11 = inst0_p15;
assign p25 = inst0_p29;
assign p5 = inst0_p9;
assign p36 = inst0_p40;
assign p8 = inst0_p12;
assign p10 = inst0_p14;
assign p7 = inst0_p11;
assign p13 = inst0_p17;
assign p18 = inst0_p22;
assign p30 = inst0_p34;
assign p24 = inst0_p28;
assign p32 = inst0_p36;
assign p14 = inst0_p18;
assign p26 = inst0_p30;
assign p31 = inst0_p35;
assign p27 = inst0_p31;
assign p33 = inst0_p37;
assign p22 = inst0_p26;
assign p34 = inst0_p38;
assign p35 = inst0_p39;
assign inst0_clk = clk;
assign inst0_p8 = p4;
assign inst0_reset = reset;
// COMPONENT END: comp93
endmodule
module comp35(
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  input logic ev0,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp35
logic ev00__0;
logic ev00__1;
logic ev00__2;
logic ev00__3;
logic ev00__4;
logic ev00_clk;
logic ev00_reset;
logic ev00_go;
logic ev00_done;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic inst1_clk;
logic inst1_reset;
fsm_5 ev00 (
    ._0(ev00__0),
    ._1(ev00__1),
    ._2(ev00__2),
    ._3(ev00__3),
    ._4(ev00__4),
    .clk(ev00_clk),
    .done(ev00_done),
    .go(ev00_go),
    .reset(ev00_reset)
);
comp34 inst1 (
    .clk(inst1_clk),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .reset(inst1_reset)
);
wire _guard0 = 1;
wire _guard1 = ev00__4;
wire _guard2 = ev00__4;
wire _guard3 = ev00__4;
wire _guard4 = ev00__4;
wire _guard5 = ev00__0;
wire _guard6 = ev00__0;
wire _guard7 = ev00__0;
wire _guard8 = ev00__0;
wire _guard9 = ev00__0;
wire _guard10 = ev00__0;
assign p16 =
  _guard1 ? inst1_p28 :
  32'd0;
assign p15 =
  _guard2 ? inst1_p27 :
  32'd0;
assign p17 =
  _guard3 ? inst1_p29 :
  32'd0;
assign p14 =
  _guard4 ? inst1_p26 :
  32'd0;
assign inst1_p20 = p8;
assign inst1_p21 = p9;
assign inst1_p23 = p11;
assign inst1_clk = clk;
assign inst1_p25 = p13;
assign inst1_reset = reset;
assign inst1_p24 = p12;
assign inst1_p22 = p10;
assign ev00_clk = clk;
assign ev00_go = ev0;
assign ev00_reset = reset;
// COMPONENT END: comp35
endmodule
module comp92(
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  output logic [1023:0] p37,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp92
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [31:0] inst0_p38;
logic [1023:0] inst0_p39;
logic inst0_clk;
logic inst0_reset;
comp91 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p39(inst0_p39),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
wire _guard0 = 1;
assign p37 = inst0_p39;
assign inst0_p19 = p17;
assign inst0_p28 = p26;
assign inst0_p29 = p27;
assign inst0_p38 = p36;
assign inst0_p12 = p10;
assign inst0_p16 = p14;
assign inst0_p9 = p7;
assign inst0_p15 = p13;
assign inst0_p17 = p15;
assign inst0_p20 = p18;
assign inst0_p21 = p19;
assign inst0_p23 = p21;
assign inst0_clk = clk;
assign inst0_p11 = p9;
assign inst0_p25 = p23;
assign inst0_p36 = p34;
assign inst0_p8 = p6;
assign inst0_p10 = p8;
assign inst0_reset = reset;
assign inst0_p7 = p5;
assign inst0_p13 = p11;
assign inst0_p18 = p16;
assign inst0_p30 = p28;
assign inst0_p24 = p22;
assign inst0_p32 = p30;
assign inst0_p14 = p12;
assign inst0_p26 = p24;
assign inst0_p31 = p29;
assign inst0_p27 = p25;
assign inst0_p33 = p31;
assign inst0_p22 = p20;
assign inst0_p34 = p32;
assign inst0_p35 = p33;
assign inst0_p37 = p35;
// COMPONENT END: comp92
endmodule
module comp57(
  input logic [127:0] p4,
  output logic [31:0] p5,
  output logic [31:0] p6,
  output logic [31:0] p7,
  output logic [31:0] p8,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp57
logic [127:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic inst0_clk;
logic inst0_reset;
comp4 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
wire _guard0 = 1;
assign p6 = inst0_p10;
assign p5 = inst0_p9;
assign p8 = inst0_p12;
assign p7 = inst0_p11;
assign inst0_clk = clk;
assign inst0_p8 = p4;
assign inst0_reset = reset;
// COMPONENT END: comp57
endmodule
module comp55(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp55
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p12;
assign p29 = p13;
assign p20 = p4;
assign p21 = p5;
assign p23 = p7;
assign p25 = p9;
assign p18 = p2;
assign p30 = p14;
assign p24 = p8;
assign p32 = p16;
assign p26 = p10;
assign p31 = p15;
assign p27 = p11;
assign p33 = p17;
assign p22 = p6;
// COMPONENT END: comp55
endmodule
module comp49(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  output logic [31:0] p40,
  output logic [31:0] p41,
  output logic [31:0] p42,
  output logic [31:0] p43,
  output logic [31:0] p44,
  output logic [31:0] p45,
  output logic [31:0] p46,
  output logic [31:0] p47,
  output logic [31:0] p48,
  output logic [31:0] p49,
  output logic [31:0] p50,
  output logic [31:0] p51,
  output logic [31:0] p52,
  output logic [31:0] p53,
  output logic [31:0] p54,
  output logic [31:0] p55,
  output logic [31:0] p56,
  output logic [31:0] p57,
  output logic [31:0] p58,
  output logic [31:0] p59,
  output logic [31:0] p60,
  output logic [31:0] p61,
  output logic [31:0] p62,
  output logic [31:0] p63,
  output logic [31:0] p64,
  output logic [31:0] p65,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp49
wire _guard0 = 1;
assign p38 = p10;
assign p40 = p14;
assign p47 = p27;
assign p65 = p33;
assign p52 = p8;
assign p59 = p21;
assign p56 = p16;
assign p60 = p24;
assign p64 = p32;
assign p36 = p6;
assign p39 = p11;
assign p46 = p26;
assign p51 = p5;
assign p54 = p12;
assign p45 = p23;
assign p53 = p9;
assign p58 = p20;
assign p50 = p4;
assign p41 = p15;
assign p43 = p19;
assign p63 = p29;
assign p42 = p18;
assign p48 = p30;
assign p49 = p31;
assign p61 = p25;
assign p62 = p28;
assign p34 = p2;
assign p35 = p3;
assign p57 = p17;
assign p37 = p7;
assign p44 = p22;
assign p55 = p13;
// COMPONENT END: comp49
endmodule
module comp63(
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  output logic [127:0] p9,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp63
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [127:0] inst0_p11;
logic inst0_clk;
logic inst0_reset;
comp62 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
wire _guard0 = 1;
assign p9 = inst0_p11;
assign inst0_p9 = p7;
assign inst0_clk = clk;
assign inst0_p8 = p6;
assign inst0_p10 = p8;
assign inst0_reset = reset;
assign inst0_p7 = p5;
// COMPONENT END: comp63
endmodule
module comp54(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp54
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p10;
assign p29 = p11;
assign p20 = p2;
assign p21 = p3;
assign p23 = p7;
assign p25 = p7;
assign p18 = p2;
assign p30 = p14;
assign p24 = p6;
assign p32 = p14;
assign p26 = p10;
assign p31 = p15;
assign p27 = p11;
assign p33 = p15;
assign p22 = p6;
// COMPONENT END: comp54
endmodule
module comp94(
  input logic [31:0] p528,
  input logic [31:0] p529,
  input logic [31:0] p530,
  input logic [31:0] p531,
  input logic [31:0] p532,
  input logic [31:0] p533,
  input logic [31:0] p534,
  input logic [31:0] p535,
  input logic [31:0] p536,
  input logic [31:0] p537,
  input logic [31:0] p538,
  input logic [31:0] p539,
  input logic [31:0] p540,
  input logic [31:0] p541,
  input logic [31:0] p542,
  input logic [31:0] p543,
  input logic [31:0] p544,
  input logic [31:0] p545,
  input logic [31:0] p546,
  input logic [31:0] p547,
  input logic [31:0] p548,
  input logic [31:0] p549,
  input logic [31:0] p550,
  input logic [31:0] p551,
  input logic [31:0] p552,
  input logic [31:0] p553,
  input logic [31:0] p554,
  input logic [31:0] p555,
  input logic [31:0] p556,
  input logic [31:0] p557,
  input logic [31:0] p558,
  input logic [31:0] p559,
  output logic [31:0] p560,
  output logic [31:0] p561,
  output logic [31:0] p562,
  output logic [31:0] p563,
  output logic [31:0] p564,
  output logic [31:0] p565,
  output logic [31:0] p566,
  output logic [31:0] p567,
  output logic [31:0] p568,
  output logic [31:0] p569,
  output logic [31:0] p570,
  output logic [31:0] p571,
  output logic [31:0] p572,
  output logic [31:0] p573,
  output logic [31:0] p574,
  output logic [31:0] p575,
  output logic [31:0] p576,
  output logic [31:0] p577,
  output logic [31:0] p578,
  output logic [31:0] p579,
  output logic [31:0] p580,
  output logic [31:0] p581,
  output logic [31:0] p582,
  output logic [31:0] p583,
  output logic [31:0] p584,
  output logic [31:0] p585,
  output logic [31:0] p586,
  output logic [31:0] p587,
  output logic [31:0] p588,
  output logic [31:0] p589,
  output logic [31:0] p590,
  output logic [31:0] p591,
  input logic ev0,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp94
logic [5:0] ev00__0state;
logic ev00__0_0;
logic [5:0] ev00__1state;
logic ev00__1_0;
logic ev00_clk;
logic ev00_reset;
logic ev00_go;
logic ev00_done;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic inst0_ev0;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_p17;
logic [31:0] inst1_p18;
logic [31:0] inst1_p19;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic [31:0] inst1_p30;
logic [31:0] inst1_p31;
logic [31:0] inst1_p32;
logic inst1_clk;
logic inst1_reset;
logic [31:0] inst2_p2;
logic [31:0] inst2_p3;
logic [31:0] inst2_p4;
logic [31:0] inst2_p5;
logic [31:0] inst2_p6;
logic [31:0] inst2_p7;
logic [31:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic [31:0] inst2_p38;
logic [31:0] inst2_p39;
logic [31:0] inst2_p40;
logic [31:0] inst2_p41;
logic [31:0] inst2_p42;
logic [31:0] inst2_p43;
logic [31:0] inst2_p44;
logic [31:0] inst2_p45;
logic [31:0] inst2_p46;
logic [31:0] inst2_p47;
logic [31:0] inst2_p48;
logic [31:0] inst2_p49;
logic [31:0] inst2_p50;
logic [31:0] inst2_p51;
logic [31:0] inst2_p52;
logic [31:0] inst2_p53;
logic [31:0] inst2_p54;
logic [31:0] inst2_p55;
logic [31:0] inst2_p56;
logic [31:0] inst2_p57;
logic [31:0] inst2_p58;
logic [31:0] inst2_p59;
logic [31:0] inst2_p60;
logic [31:0] inst2_p61;
logic [31:0] inst2_p62;
logic [31:0] inst2_p63;
logic [31:0] inst2_p64;
logic [31:0] inst2_p65;
logic inst2_clk;
logic inst2_reset;
logic [31:0] inst3_p2;
logic [31:0] inst3_p3;
logic [31:0] inst3_p4;
logic [31:0] inst3_p5;
logic [31:0] inst3_p6;
logic [31:0] inst3_p7;
logic [31:0] inst3_p8;
logic [31:0] inst3_p9;
logic [31:0] inst3_p10;
logic [31:0] inst3_p11;
logic [31:0] inst3_p12;
logic [31:0] inst3_p13;
logic [31:0] inst3_p14;
logic [31:0] inst3_p15;
logic [31:0] inst3_p16;
logic [31:0] inst3_p17;
logic [31:0] inst3_p18;
logic [31:0] inst3_p19;
logic [31:0] inst3_p20;
logic [31:0] inst3_p21;
logic [31:0] inst3_p22;
logic [31:0] inst3_p23;
logic [31:0] inst3_p24;
logic [31:0] inst3_p25;
logic [31:0] inst3_p26;
logic [31:0] inst3_p27;
logic [31:0] inst3_p28;
logic [31:0] inst3_p29;
logic [31:0] inst3_p30;
logic [31:0] inst3_p31;
logic [31:0] inst3_p32;
logic [31:0] inst3_p33;
logic [31:0] inst3_p34;
logic [31:0] inst3_p35;
logic [31:0] inst3_p36;
logic [31:0] inst3_p37;
logic [31:0] inst3_p38;
logic [31:0] inst3_p39;
logic [31:0] inst3_p40;
logic [31:0] inst3_p41;
logic [31:0] inst3_p42;
logic [31:0] inst3_p43;
logic [31:0] inst3_p44;
logic [31:0] inst3_p45;
logic [31:0] inst3_p46;
logic [31:0] inst3_p47;
logic [31:0] inst3_p48;
logic [31:0] inst3_p49;
logic [31:0] inst3_p50;
logic [31:0] inst3_p51;
logic [31:0] inst3_p52;
logic [31:0] inst3_p53;
logic [31:0] inst3_p54;
logic [31:0] inst3_p55;
logic [31:0] inst3_p56;
logic [31:0] inst3_p57;
logic [31:0] inst3_p58;
logic [31:0] inst3_p59;
logic [31:0] inst3_p60;
logic [31:0] inst3_p61;
logic [31:0] inst3_p62;
logic [31:0] inst3_p63;
logic [31:0] inst3_p64;
logic [31:0] inst3_p65;
logic inst3_reset;
logic inst3_clk;
logic [1023:0] inst4_in;
logic [1023:0] inst4_out;
logic inst4_clk;
logic inst4_reset;
logic [31:0] inst5_p2;
logic [31:0] inst5_p3;
logic [31:0] inst5_p4;
logic [31:0] inst5_p5;
logic [31:0] inst5_p6;
logic [31:0] inst5_p7;
logic [31:0] inst5_p8;
logic [31:0] inst5_p9;
logic [31:0] inst5_p10;
logic [31:0] inst5_p11;
logic [31:0] inst5_p12;
logic [31:0] inst5_p13;
logic [31:0] inst5_p14;
logic [31:0] inst5_p15;
logic [31:0] inst5_p16;
logic [31:0] inst5_p17;
logic [31:0] inst5_p18;
logic [31:0] inst5_p19;
logic [31:0] inst5_p20;
logic [31:0] inst5_p21;
logic [31:0] inst5_p22;
logic [31:0] inst5_p23;
logic [31:0] inst5_p24;
logic [31:0] inst5_p25;
logic [31:0] inst5_p26;
logic [31:0] inst5_p27;
logic [31:0] inst5_p28;
logic [31:0] inst5_p29;
logic [31:0] inst5_p30;
logic [31:0] inst5_p31;
logic [31:0] inst5_p32;
logic [31:0] inst5_p33;
logic inst5_reset;
logic inst5_clk;
logic [31:0] inst6_p2;
logic [31:0] inst6_p3;
logic [31:0] inst6_p4;
logic [31:0] inst6_p5;
logic [31:0] inst6_p6;
logic [31:0] inst6_p7;
logic [31:0] inst6_p8;
logic [31:0] inst6_p9;
logic [31:0] inst6_p10;
logic [31:0] inst6_p11;
logic [31:0] inst6_p12;
logic [31:0] inst6_p13;
logic [31:0] inst6_p14;
logic [31:0] inst6_p15;
logic [31:0] inst6_p16;
logic [31:0] inst6_p17;
logic [31:0] inst6_p18;
logic [31:0] inst6_p19;
logic [31:0] inst6_p20;
logic [31:0] inst6_p21;
logic [31:0] inst6_p22;
logic [31:0] inst6_p23;
logic [31:0] inst6_p24;
logic [31:0] inst6_p25;
logic [31:0] inst6_p26;
logic [31:0] inst6_p27;
logic [31:0] inst6_p28;
logic [31:0] inst6_p29;
logic [31:0] inst6_p30;
logic [31:0] inst6_p31;
logic [31:0] inst6_p32;
logic [31:0] inst6_p33;
logic inst6_clk;
logic inst6_reset;
logic [31:0] inst7_p2;
logic [31:0] inst7_p3;
logic [31:0] inst7_p4;
logic [31:0] inst7_p5;
logic [31:0] inst7_p6;
logic [31:0] inst7_p7;
logic [31:0] inst7_p8;
logic [31:0] inst7_p9;
logic [31:0] inst7_p10;
logic [31:0] inst7_p11;
logic [31:0] inst7_p12;
logic [31:0] inst7_p13;
logic [31:0] inst7_p14;
logic [31:0] inst7_p15;
logic [31:0] inst7_p16;
logic [31:0] inst7_p17;
logic [31:0] inst7_p18;
logic [31:0] inst7_p19;
logic [31:0] inst7_p20;
logic [31:0] inst7_p21;
logic [31:0] inst7_p22;
logic [31:0] inst7_p23;
logic [31:0] inst7_p24;
logic [31:0] inst7_p25;
logic [31:0] inst7_p26;
logic [31:0] inst7_p27;
logic [31:0] inst7_p28;
logic [31:0] inst7_p29;
logic [31:0] inst7_p30;
logic [31:0] inst7_p31;
logic [31:0] inst7_p32;
logic [31:0] inst7_p33;
logic inst7_clk;
logic inst7_reset;
logic [31:0] inst8_p2;
logic [31:0] inst8_p3;
logic [31:0] inst8_p4;
logic [31:0] inst8_p5;
logic [31:0] inst8_p6;
logic [31:0] inst8_p7;
logic [31:0] inst8_p8;
logic [31:0] inst8_p9;
logic [31:0] inst8_p10;
logic [31:0] inst8_p11;
logic [31:0] inst8_p12;
logic [31:0] inst8_p13;
logic [31:0] inst8_p14;
logic [31:0] inst8_p15;
logic [31:0] inst8_p16;
logic [31:0] inst8_p17;
logic [31:0] inst8_p18;
logic [31:0] inst8_p19;
logic [31:0] inst8_p20;
logic [31:0] inst8_p21;
logic [31:0] inst8_p22;
logic [31:0] inst8_p23;
logic [31:0] inst8_p24;
logic [31:0] inst8_p25;
logic [31:0] inst8_p26;
logic [31:0] inst8_p27;
logic [31:0] inst8_p28;
logic [31:0] inst8_p29;
logic [31:0] inst8_p30;
logic [31:0] inst8_p31;
logic [31:0] inst8_p32;
logic [31:0] inst8_p33;
logic inst8_clk;
logic inst8_reset;
logic [127:0] inst9_in;
logic [127:0] inst9_out;
logic inst9_clk;
logic inst9_reset;
logic inst9_write_en;
logic [127:0] inst10_p4;
logic [31:0] inst10_p5;
logic [31:0] inst10_p6;
logic [31:0] inst10_p7;
logic [31:0] inst10_p8;
logic inst10_reset;
logic inst10_clk;
logic [31:0] inst11_p5;
logic [31:0] inst11_p6;
logic [31:0] inst11_p7;
logic [31:0] inst11_p8;
logic [127:0] inst11_p9;
logic inst11_clk;
logic inst11_reset;
logic [31:0] inst12_p5;
logic [31:0] inst12_p6;
logic [31:0] inst12_p7;
logic [31:0] inst12_p8;
logic [127:0] inst12_p9;
logic inst12_clk;
logic inst12_reset;
logic [127:0] inst13_p4;
logic [31:0] inst13_p5;
logic [31:0] inst13_p6;
logic [31:0] inst13_p7;
logic [31:0] inst13_p8;
logic inst13_reset;
logic inst13_clk;
logic [127:0] inst14_p4;
logic [31:0] inst14_p5;
logic [31:0] inst14_p6;
logic [31:0] inst14_p7;
logic [31:0] inst14_p8;
logic inst14_reset;
logic inst14_clk;
logic [31:0] inst15_p5;
logic [31:0] inst15_p6;
logic [31:0] inst15_p7;
logic [31:0] inst15_p8;
logic [127:0] inst15_p9;
logic inst15_clk;
logic inst15_reset;
logic [31:0] inst16_p5;
logic [31:0] inst16_p6;
logic [31:0] inst16_p7;
logic [31:0] inst16_p8;
logic [127:0] inst16_p9;
logic inst16_clk;
logic inst16_reset;
logic [127:0] inst17_p4;
logic [31:0] inst17_p5;
logic [31:0] inst17_p6;
logic [31:0] inst17_p7;
logic [31:0] inst17_p8;
logic inst17_reset;
logic inst17_clk;
logic [127:0] inst18_p4;
logic [31:0] inst18_p5;
logic [31:0] inst18_p6;
logic [31:0] inst18_p7;
logic [31:0] inst18_p8;
logic inst18_reset;
logic inst18_clk;
logic [31:0] inst19_p5;
logic [31:0] inst19_p6;
logic [31:0] inst19_p7;
logic [31:0] inst19_p8;
logic [127:0] inst19_p9;
logic inst19_clk;
logic inst19_reset;
logic [31:0] inst20_p5;
logic [31:0] inst20_p6;
logic [31:0] inst20_p7;
logic [31:0] inst20_p8;
logic [127:0] inst20_p9;
logic inst20_clk;
logic inst20_reset;
logic [127:0] inst21_p4;
logic [31:0] inst21_p5;
logic [31:0] inst21_p6;
logic [31:0] inst21_p7;
logic [31:0] inst21_p8;
logic inst21_reset;
logic inst21_clk;
logic [127:0] inst22_p4;
logic [31:0] inst22_p5;
logic [31:0] inst22_p6;
logic [31:0] inst22_p7;
logic [31:0] inst22_p8;
logic inst22_reset;
logic inst22_clk;
logic [31:0] inst23_p5;
logic [31:0] inst23_p6;
logic [31:0] inst23_p7;
logic [31:0] inst23_p8;
logic [127:0] inst23_p9;
logic inst23_clk;
logic inst23_reset;
logic [31:0] inst24_p5;
logic [31:0] inst24_p6;
logic [31:0] inst24_p7;
logic [31:0] inst24_p8;
logic [127:0] inst24_p9;
logic inst24_clk;
logic inst24_reset;
logic [127:0] inst25_p4;
logic [31:0] inst25_p5;
logic [31:0] inst25_p6;
logic [31:0] inst25_p7;
logic [31:0] inst25_p8;
logic inst25_reset;
logic inst25_clk;
logic [127:0] inst26_in;
logic [127:0] inst26_out;
logic inst26_clk;
logic inst26_reset;
logic inst26_write_en;
logic [127:0] inst27_p4;
logic [31:0] inst27_p5;
logic [31:0] inst27_p6;
logic [31:0] inst27_p7;
logic [31:0] inst27_p8;
logic inst27_reset;
logic inst27_clk;
logic [31:0] inst28_p5;
logic [31:0] inst28_p6;
logic [31:0] inst28_p7;
logic [31:0] inst28_p8;
logic [127:0] inst28_p9;
logic inst28_clk;
logic inst28_reset;
logic [31:0] inst29_p5;
logic [31:0] inst29_p6;
logic [31:0] inst29_p7;
logic [31:0] inst29_p8;
logic [127:0] inst29_p9;
logic inst29_clk;
logic inst29_reset;
logic [127:0] inst30_p4;
logic [31:0] inst30_p5;
logic [31:0] inst30_p6;
logic [31:0] inst30_p7;
logic [31:0] inst30_p8;
logic inst30_reset;
logic inst30_clk;
logic [127:0] inst31_p4;
logic [31:0] inst31_p5;
logic [31:0] inst31_p6;
logic [31:0] inst31_p7;
logic [31:0] inst31_p8;
logic inst31_reset;
logic inst31_clk;
logic [31:0] inst32_p5;
logic [31:0] inst32_p6;
logic [31:0] inst32_p7;
logic [31:0] inst32_p8;
logic [127:0] inst32_p9;
logic inst32_clk;
logic inst32_reset;
logic [31:0] inst33_p5;
logic [31:0] inst33_p6;
logic [31:0] inst33_p7;
logic [31:0] inst33_p8;
logic [127:0] inst33_p9;
logic inst33_clk;
logic inst33_reset;
logic [127:0] inst34_p4;
logic [31:0] inst34_p5;
logic [31:0] inst34_p6;
logic [31:0] inst34_p7;
logic [31:0] inst34_p8;
logic inst34_reset;
logic inst34_clk;
logic [127:0] inst35_p4;
logic [31:0] inst35_p5;
logic [31:0] inst35_p6;
logic [31:0] inst35_p7;
logic [31:0] inst35_p8;
logic inst35_reset;
logic inst35_clk;
logic [31:0] inst36_p5;
logic [31:0] inst36_p6;
logic [31:0] inst36_p7;
logic [31:0] inst36_p8;
logic [127:0] inst36_p9;
logic inst36_clk;
logic inst36_reset;
logic [31:0] inst37_p5;
logic [31:0] inst37_p6;
logic [31:0] inst37_p7;
logic [31:0] inst37_p8;
logic [127:0] inst37_p9;
logic inst37_clk;
logic inst37_reset;
logic [127:0] inst38_p4;
logic [31:0] inst38_p5;
logic [31:0] inst38_p6;
logic [31:0] inst38_p7;
logic [31:0] inst38_p8;
logic inst38_reset;
logic inst38_clk;
logic [127:0] inst39_p4;
logic [31:0] inst39_p5;
logic [31:0] inst39_p6;
logic [31:0] inst39_p7;
logic [31:0] inst39_p8;
logic inst39_reset;
logic inst39_clk;
logic [31:0] inst40_p5;
logic [31:0] inst40_p6;
logic [31:0] inst40_p7;
logic [31:0] inst40_p8;
logic [127:0] inst40_p9;
logic inst40_clk;
logic inst40_reset;
logic [31:0] inst41_p5;
logic [31:0] inst41_p6;
logic [31:0] inst41_p7;
logic [31:0] inst41_p8;
logic [127:0] inst41_p9;
logic inst41_clk;
logic inst41_reset;
logic [127:0] inst42_p4;
logic [31:0] inst42_p5;
logic [31:0] inst42_p6;
logic [31:0] inst42_p7;
logic [31:0] inst42_p8;
logic inst42_reset;
logic inst42_clk;
logic [127:0] inst43_in;
logic [127:0] inst43_out;
logic inst43_clk;
logic inst43_reset;
logic inst43_write_en;
logic [127:0] inst44_p4;
logic [31:0] inst44_p5;
logic [31:0] inst44_p6;
logic [31:0] inst44_p7;
logic [31:0] inst44_p8;
logic inst44_reset;
logic inst44_clk;
logic [31:0] inst45_p5;
logic [31:0] inst45_p6;
logic [31:0] inst45_p7;
logic [31:0] inst45_p8;
logic [127:0] inst45_p9;
logic inst45_clk;
logic inst45_reset;
logic [31:0] inst46_p5;
logic [31:0] inst46_p6;
logic [31:0] inst46_p7;
logic [31:0] inst46_p8;
logic [127:0] inst46_p9;
logic inst46_clk;
logic inst46_reset;
logic [127:0] inst47_p4;
logic [31:0] inst47_p5;
logic [31:0] inst47_p6;
logic [31:0] inst47_p7;
logic [31:0] inst47_p8;
logic inst47_reset;
logic inst47_clk;
logic [127:0] inst48_p4;
logic [31:0] inst48_p5;
logic [31:0] inst48_p6;
logic [31:0] inst48_p7;
logic [31:0] inst48_p8;
logic inst48_reset;
logic inst48_clk;
logic [31:0] inst49_p5;
logic [31:0] inst49_p6;
logic [31:0] inst49_p7;
logic [31:0] inst49_p8;
logic [127:0] inst49_p9;
logic inst49_clk;
logic inst49_reset;
logic [31:0] inst50_p5;
logic [31:0] inst50_p6;
logic [31:0] inst50_p7;
logic [31:0] inst50_p8;
logic [127:0] inst50_p9;
logic inst50_clk;
logic inst50_reset;
logic [127:0] inst51_p4;
logic [31:0] inst51_p5;
logic [31:0] inst51_p6;
logic [31:0] inst51_p7;
logic [31:0] inst51_p8;
logic inst51_reset;
logic inst51_clk;
logic [127:0] inst52_p4;
logic [31:0] inst52_p5;
logic [31:0] inst52_p6;
logic [31:0] inst52_p7;
logic [31:0] inst52_p8;
logic inst52_reset;
logic inst52_clk;
logic [31:0] inst53_p5;
logic [31:0] inst53_p6;
logic [31:0] inst53_p7;
logic [31:0] inst53_p8;
logic [127:0] inst53_p9;
logic inst53_clk;
logic inst53_reset;
logic [31:0] inst54_p5;
logic [31:0] inst54_p6;
logic [31:0] inst54_p7;
logic [31:0] inst54_p8;
logic [127:0] inst54_p9;
logic inst54_clk;
logic inst54_reset;
logic [127:0] inst55_p4;
logic [31:0] inst55_p5;
logic [31:0] inst55_p6;
logic [31:0] inst55_p7;
logic [31:0] inst55_p8;
logic inst55_reset;
logic inst55_clk;
logic [127:0] inst56_p4;
logic [31:0] inst56_p5;
logic [31:0] inst56_p6;
logic [31:0] inst56_p7;
logic [31:0] inst56_p8;
logic inst56_reset;
logic inst56_clk;
logic [31:0] inst57_p5;
logic [31:0] inst57_p6;
logic [31:0] inst57_p7;
logic [31:0] inst57_p8;
logic [127:0] inst57_p9;
logic inst57_clk;
logic inst57_reset;
logic [31:0] inst58_p5;
logic [31:0] inst58_p6;
logic [31:0] inst58_p7;
logic [31:0] inst58_p8;
logic [127:0] inst58_p9;
logic inst58_clk;
logic inst58_reset;
logic [127:0] inst59_p4;
logic [31:0] inst59_p5;
logic [31:0] inst59_p6;
logic [31:0] inst59_p7;
logic [31:0] inst59_p8;
logic inst59_reset;
logic inst59_clk;
logic [127:0] inst60_in;
logic [127:0] inst60_out;
logic inst60_clk;
logic inst60_reset;
logic inst60_write_en;
logic [127:0] inst61_p4;
logic [31:0] inst61_p5;
logic [31:0] inst61_p6;
logic [31:0] inst61_p7;
logic [31:0] inst61_p8;
logic inst61_reset;
logic inst61_clk;
logic [31:0] inst62_p5;
logic [31:0] inst62_p6;
logic [31:0] inst62_p7;
logic [31:0] inst62_p8;
logic [127:0] inst62_p9;
logic inst62_clk;
logic inst62_reset;
logic [31:0] inst63_p5;
logic [31:0] inst63_p6;
logic [31:0] inst63_p7;
logic [31:0] inst63_p8;
logic [127:0] inst63_p9;
logic inst63_clk;
logic inst63_reset;
logic [127:0] inst64_p4;
logic [31:0] inst64_p5;
logic [31:0] inst64_p6;
logic [31:0] inst64_p7;
logic [31:0] inst64_p8;
logic inst64_reset;
logic inst64_clk;
logic [127:0] inst65_p4;
logic [31:0] inst65_p5;
logic [31:0] inst65_p6;
logic [31:0] inst65_p7;
logic [31:0] inst65_p8;
logic inst65_reset;
logic inst65_clk;
logic [31:0] inst66_p5;
logic [31:0] inst66_p6;
logic [31:0] inst66_p7;
logic [31:0] inst66_p8;
logic [127:0] inst66_p9;
logic inst66_clk;
logic inst66_reset;
logic [31:0] inst67_p5;
logic [31:0] inst67_p6;
logic [31:0] inst67_p7;
logic [31:0] inst67_p8;
logic [127:0] inst67_p9;
logic inst67_clk;
logic inst67_reset;
logic [127:0] inst68_p4;
logic [31:0] inst68_p5;
logic [31:0] inst68_p6;
logic [31:0] inst68_p7;
logic [31:0] inst68_p8;
logic inst68_reset;
logic inst68_clk;
logic [127:0] inst69_p4;
logic [31:0] inst69_p5;
logic [31:0] inst69_p6;
logic [31:0] inst69_p7;
logic [31:0] inst69_p8;
logic inst69_reset;
logic inst69_clk;
logic [31:0] inst70_p5;
logic [31:0] inst70_p6;
logic [31:0] inst70_p7;
logic [31:0] inst70_p8;
logic [127:0] inst70_p9;
logic inst70_clk;
logic inst70_reset;
logic [31:0] inst71_p5;
logic [31:0] inst71_p6;
logic [31:0] inst71_p7;
logic [31:0] inst71_p8;
logic [127:0] inst71_p9;
logic inst71_clk;
logic inst71_reset;
logic [127:0] inst72_p4;
logic [31:0] inst72_p5;
logic [31:0] inst72_p6;
logic [31:0] inst72_p7;
logic [31:0] inst72_p8;
logic inst72_reset;
logic inst72_clk;
logic [127:0] inst73_p4;
logic [31:0] inst73_p5;
logic [31:0] inst73_p6;
logic [31:0] inst73_p7;
logic [31:0] inst73_p8;
logic inst73_reset;
logic inst73_clk;
logic [31:0] inst74_p5;
logic [31:0] inst74_p6;
logic [31:0] inst74_p7;
logic [31:0] inst74_p8;
logic [127:0] inst74_p9;
logic inst74_clk;
logic inst74_reset;
logic [31:0] inst75_p5;
logic [31:0] inst75_p6;
logic [31:0] inst75_p7;
logic [31:0] inst75_p8;
logic [127:0] inst75_p9;
logic inst75_clk;
logic inst75_reset;
logic [127:0] inst76_p4;
logic [31:0] inst76_p5;
logic [31:0] inst76_p6;
logic [31:0] inst76_p7;
logic [31:0] inst76_p8;
logic inst76_reset;
logic inst76_clk;
logic [127:0] inst77_in;
logic [127:0] inst77_out;
logic inst77_clk;
logic inst77_reset;
logic inst77_write_en;
logic [127:0] inst78_p4;
logic [31:0] inst78_p5;
logic [31:0] inst78_p6;
logic [31:0] inst78_p7;
logic [31:0] inst78_p8;
logic inst78_reset;
logic inst78_clk;
logic [31:0] inst79_p5;
logic [31:0] inst79_p6;
logic [31:0] inst79_p7;
logic [31:0] inst79_p8;
logic [127:0] inst79_p9;
logic inst79_clk;
logic inst79_reset;
logic [31:0] inst80_p5;
logic [31:0] inst80_p6;
logic [31:0] inst80_p7;
logic [31:0] inst80_p8;
logic [127:0] inst80_p9;
logic inst80_clk;
logic inst80_reset;
logic [127:0] inst81_p4;
logic [31:0] inst81_p5;
logic [31:0] inst81_p6;
logic [31:0] inst81_p7;
logic [31:0] inst81_p8;
logic inst81_reset;
logic inst81_clk;
logic [127:0] inst82_p4;
logic [31:0] inst82_p5;
logic [31:0] inst82_p6;
logic [31:0] inst82_p7;
logic [31:0] inst82_p8;
logic inst82_reset;
logic inst82_clk;
logic [31:0] inst83_p5;
logic [31:0] inst83_p6;
logic [31:0] inst83_p7;
logic [31:0] inst83_p8;
logic [127:0] inst83_p9;
logic inst83_clk;
logic inst83_reset;
logic [31:0] inst84_p5;
logic [31:0] inst84_p6;
logic [31:0] inst84_p7;
logic [31:0] inst84_p8;
logic [127:0] inst84_p9;
logic inst84_clk;
logic inst84_reset;
logic [127:0] inst85_p4;
logic [31:0] inst85_p5;
logic [31:0] inst85_p6;
logic [31:0] inst85_p7;
logic [31:0] inst85_p8;
logic inst85_reset;
logic inst85_clk;
logic [127:0] inst86_p4;
logic [31:0] inst86_p5;
logic [31:0] inst86_p6;
logic [31:0] inst86_p7;
logic [31:0] inst86_p8;
logic inst86_reset;
logic inst86_clk;
logic [31:0] inst87_p5;
logic [31:0] inst87_p6;
logic [31:0] inst87_p7;
logic [31:0] inst87_p8;
logic [127:0] inst87_p9;
logic inst87_clk;
logic inst87_reset;
logic [31:0] inst88_p5;
logic [31:0] inst88_p6;
logic [31:0] inst88_p7;
logic [31:0] inst88_p8;
logic [127:0] inst88_p9;
logic inst88_clk;
logic inst88_reset;
logic [127:0] inst89_p4;
logic [31:0] inst89_p5;
logic [31:0] inst89_p6;
logic [31:0] inst89_p7;
logic [31:0] inst89_p8;
logic inst89_reset;
logic inst89_clk;
logic [127:0] inst90_p4;
logic [31:0] inst90_p5;
logic [31:0] inst90_p6;
logic [31:0] inst90_p7;
logic [31:0] inst90_p8;
logic inst90_reset;
logic inst90_clk;
logic [31:0] inst91_p5;
logic [31:0] inst91_p6;
logic [31:0] inst91_p7;
logic [31:0] inst91_p8;
logic [127:0] inst91_p9;
logic inst91_clk;
logic inst91_reset;
logic [31:0] inst92_p5;
logic [31:0] inst92_p6;
logic [31:0] inst92_p7;
logic [31:0] inst92_p8;
logic [127:0] inst92_p9;
logic inst92_clk;
logic inst92_reset;
logic [127:0] inst93_p4;
logic [31:0] inst93_p5;
logic [31:0] inst93_p6;
logic [31:0] inst93_p7;
logic [31:0] inst93_p8;
logic inst93_reset;
logic inst93_clk;
logic [127:0] inst94_in;
logic [127:0] inst94_out;
logic inst94_clk;
logic inst94_reset;
logic inst94_write_en;
logic [127:0] inst95_p4;
logic [31:0] inst95_p5;
logic [31:0] inst95_p6;
logic [31:0] inst95_p7;
logic [31:0] inst95_p8;
logic inst95_reset;
logic inst95_clk;
logic [31:0] inst96_p5;
logic [31:0] inst96_p6;
logic [31:0] inst96_p7;
logic [31:0] inst96_p8;
logic [127:0] inst96_p9;
logic inst96_clk;
logic inst96_reset;
logic [31:0] inst97_p5;
logic [31:0] inst97_p6;
logic [31:0] inst97_p7;
logic [31:0] inst97_p8;
logic [127:0] inst97_p9;
logic inst97_clk;
logic inst97_reset;
logic [127:0] inst98_p4;
logic [31:0] inst98_p5;
logic [31:0] inst98_p6;
logic [31:0] inst98_p7;
logic [31:0] inst98_p8;
logic inst98_reset;
logic inst98_clk;
logic [127:0] inst99_p4;
logic [31:0] inst99_p5;
logic [31:0] inst99_p6;
logic [31:0] inst99_p7;
logic [31:0] inst99_p8;
logic inst99_reset;
logic inst99_clk;
logic [31:0] inst100_p5;
logic [31:0] inst100_p6;
logic [31:0] inst100_p7;
logic [31:0] inst100_p8;
logic [127:0] inst100_p9;
logic inst100_clk;
logic inst100_reset;
logic [31:0] inst101_p5;
logic [31:0] inst101_p6;
logic [31:0] inst101_p7;
logic [31:0] inst101_p8;
logic [127:0] inst101_p9;
logic inst101_clk;
logic inst101_reset;
logic [127:0] inst102_p4;
logic [31:0] inst102_p5;
logic [31:0] inst102_p6;
logic [31:0] inst102_p7;
logic [31:0] inst102_p8;
logic inst102_reset;
logic inst102_clk;
logic [127:0] inst103_p4;
logic [31:0] inst103_p5;
logic [31:0] inst103_p6;
logic [31:0] inst103_p7;
logic [31:0] inst103_p8;
logic inst103_reset;
logic inst103_clk;
logic [31:0] inst104_p5;
logic [31:0] inst104_p6;
logic [31:0] inst104_p7;
logic [31:0] inst104_p8;
logic [127:0] inst104_p9;
logic inst104_clk;
logic inst104_reset;
logic [31:0] inst105_p5;
logic [31:0] inst105_p6;
logic [31:0] inst105_p7;
logic [31:0] inst105_p8;
logic [127:0] inst105_p9;
logic inst105_clk;
logic inst105_reset;
logic [127:0] inst106_p4;
logic [31:0] inst106_p5;
logic [31:0] inst106_p6;
logic [31:0] inst106_p7;
logic [31:0] inst106_p8;
logic inst106_reset;
logic inst106_clk;
logic [127:0] inst107_p4;
logic [31:0] inst107_p5;
logic [31:0] inst107_p6;
logic [31:0] inst107_p7;
logic [31:0] inst107_p8;
logic inst107_reset;
logic inst107_clk;
logic [31:0] inst108_p5;
logic [31:0] inst108_p6;
logic [31:0] inst108_p7;
logic [31:0] inst108_p8;
logic [127:0] inst108_p9;
logic inst108_clk;
logic inst108_reset;
logic [31:0] inst109_p5;
logic [31:0] inst109_p6;
logic [31:0] inst109_p7;
logic [31:0] inst109_p8;
logic [127:0] inst109_p9;
logic inst109_clk;
logic inst109_reset;
logic [127:0] inst110_p4;
logic [31:0] inst110_p5;
logic [31:0] inst110_p6;
logic [31:0] inst110_p7;
logic [31:0] inst110_p8;
logic inst110_reset;
logic inst110_clk;
logic [127:0] inst111_in;
logic [127:0] inst111_out;
logic inst111_clk;
logic inst111_reset;
logic inst111_write_en;
logic [127:0] inst112_p4;
logic [31:0] inst112_p5;
logic [31:0] inst112_p6;
logic [31:0] inst112_p7;
logic [31:0] inst112_p8;
logic inst112_reset;
logic inst112_clk;
logic [31:0] inst113_p5;
logic [31:0] inst113_p6;
logic [31:0] inst113_p7;
logic [31:0] inst113_p8;
logic [127:0] inst113_p9;
logic inst113_clk;
logic inst113_reset;
logic [31:0] inst114_p5;
logic [31:0] inst114_p6;
logic [31:0] inst114_p7;
logic [31:0] inst114_p8;
logic [127:0] inst114_p9;
logic inst114_clk;
logic inst114_reset;
logic [127:0] inst115_p4;
logic [31:0] inst115_p5;
logic [31:0] inst115_p6;
logic [31:0] inst115_p7;
logic [31:0] inst115_p8;
logic inst115_reset;
logic inst115_clk;
logic [127:0] inst116_p4;
logic [31:0] inst116_p5;
logic [31:0] inst116_p6;
logic [31:0] inst116_p7;
logic [31:0] inst116_p8;
logic inst116_reset;
logic inst116_clk;
logic [31:0] inst117_p5;
logic [31:0] inst117_p6;
logic [31:0] inst117_p7;
logic [31:0] inst117_p8;
logic [127:0] inst117_p9;
logic inst117_clk;
logic inst117_reset;
logic [31:0] inst118_p5;
logic [31:0] inst118_p6;
logic [31:0] inst118_p7;
logic [31:0] inst118_p8;
logic [127:0] inst118_p9;
logic inst118_clk;
logic inst118_reset;
logic [127:0] inst119_p4;
logic [31:0] inst119_p5;
logic [31:0] inst119_p6;
logic [31:0] inst119_p7;
logic [31:0] inst119_p8;
logic inst119_reset;
logic inst119_clk;
logic [127:0] inst120_p4;
logic [31:0] inst120_p5;
logic [31:0] inst120_p6;
logic [31:0] inst120_p7;
logic [31:0] inst120_p8;
logic inst120_reset;
logic inst120_clk;
logic [31:0] inst121_p5;
logic [31:0] inst121_p6;
logic [31:0] inst121_p7;
logic [31:0] inst121_p8;
logic [127:0] inst121_p9;
logic inst121_clk;
logic inst121_reset;
logic [31:0] inst122_p5;
logic [31:0] inst122_p6;
logic [31:0] inst122_p7;
logic [31:0] inst122_p8;
logic [127:0] inst122_p9;
logic inst122_clk;
logic inst122_reset;
logic [127:0] inst123_p4;
logic [31:0] inst123_p5;
logic [31:0] inst123_p6;
logic [31:0] inst123_p7;
logic [31:0] inst123_p8;
logic inst123_reset;
logic inst123_clk;
logic [127:0] inst124_p4;
logic [31:0] inst124_p5;
logic [31:0] inst124_p6;
logic [31:0] inst124_p7;
logic [31:0] inst124_p8;
logic inst124_reset;
logic inst124_clk;
logic [31:0] inst125_p5;
logic [31:0] inst125_p6;
logic [31:0] inst125_p7;
logic [31:0] inst125_p8;
logic [127:0] inst125_p9;
logic inst125_clk;
logic inst125_reset;
logic [31:0] inst126_p5;
logic [31:0] inst126_p6;
logic [31:0] inst126_p7;
logic [31:0] inst126_p8;
logic [127:0] inst126_p9;
logic inst126_clk;
logic inst126_reset;
logic [127:0] inst127_p4;
logic [31:0] inst127_p5;
logic [31:0] inst127_p6;
logic [31:0] inst127_p7;
logic [31:0] inst127_p8;
logic inst127_reset;
logic inst127_clk;
logic [127:0] inst128_in;
logic [127:0] inst128_out;
logic inst128_clk;
logic inst128_reset;
logic inst128_write_en;
logic [127:0] inst129_p4;
logic [31:0] inst129_p5;
logic [31:0] inst129_p6;
logic [31:0] inst129_p7;
logic [31:0] inst129_p8;
logic inst129_reset;
logic inst129_clk;
logic [31:0] inst130_p5;
logic [31:0] inst130_p6;
logic [31:0] inst130_p7;
logic [31:0] inst130_p8;
logic [127:0] inst130_p9;
logic inst130_clk;
logic inst130_reset;
logic [31:0] inst131_p5;
logic [31:0] inst131_p6;
logic [31:0] inst131_p7;
logic [31:0] inst131_p8;
logic [127:0] inst131_p9;
logic inst131_clk;
logic inst131_reset;
logic [127:0] inst132_p4;
logic [31:0] inst132_p5;
logic [31:0] inst132_p6;
logic [31:0] inst132_p7;
logic [31:0] inst132_p8;
logic inst132_reset;
logic inst132_clk;
logic [127:0] inst133_p4;
logic [31:0] inst133_p5;
logic [31:0] inst133_p6;
logic [31:0] inst133_p7;
logic [31:0] inst133_p8;
logic inst133_reset;
logic inst133_clk;
logic [31:0] inst134_p5;
logic [31:0] inst134_p6;
logic [31:0] inst134_p7;
logic [31:0] inst134_p8;
logic [127:0] inst134_p9;
logic inst134_clk;
logic inst134_reset;
logic [31:0] inst135_p5;
logic [31:0] inst135_p6;
logic [31:0] inst135_p7;
logic [31:0] inst135_p8;
logic [127:0] inst135_p9;
logic inst135_clk;
logic inst135_reset;
logic [127:0] inst136_p4;
logic [31:0] inst136_p5;
logic [31:0] inst136_p6;
logic [31:0] inst136_p7;
logic [31:0] inst136_p8;
logic inst136_reset;
logic inst136_clk;
logic [127:0] inst137_p4;
logic [31:0] inst137_p5;
logic [31:0] inst137_p6;
logic [31:0] inst137_p7;
logic [31:0] inst137_p8;
logic inst137_reset;
logic inst137_clk;
logic [31:0] inst138_p5;
logic [31:0] inst138_p6;
logic [31:0] inst138_p7;
logic [31:0] inst138_p8;
logic [127:0] inst138_p9;
logic inst138_clk;
logic inst138_reset;
logic [31:0] inst139_p5;
logic [31:0] inst139_p6;
logic [31:0] inst139_p7;
logic [31:0] inst139_p8;
logic [127:0] inst139_p9;
logic inst139_clk;
logic inst139_reset;
logic [127:0] inst140_p4;
logic [31:0] inst140_p5;
logic [31:0] inst140_p6;
logic [31:0] inst140_p7;
logic [31:0] inst140_p8;
logic inst140_reset;
logic inst140_clk;
logic [127:0] inst141_p4;
logic [31:0] inst141_p5;
logic [31:0] inst141_p6;
logic [31:0] inst141_p7;
logic [31:0] inst141_p8;
logic inst141_reset;
logic inst141_clk;
logic [31:0] inst142_p5;
logic [31:0] inst142_p6;
logic [31:0] inst142_p7;
logic [31:0] inst142_p8;
logic [127:0] inst142_p9;
logic inst142_clk;
logic inst142_reset;
logic [31:0] inst143_p5;
logic [31:0] inst143_p6;
logic [31:0] inst143_p7;
logic [31:0] inst143_p8;
logic [127:0] inst143_p9;
logic inst143_clk;
logic inst143_reset;
logic [127:0] inst144_p4;
logic [31:0] inst144_p5;
logic [31:0] inst144_p6;
logic [31:0] inst144_p7;
logic [31:0] inst144_p8;
logic inst144_reset;
logic inst144_clk;
logic [31:0] inst145_p5;
logic [31:0] inst145_p6;
logic [31:0] inst145_p7;
logic [31:0] inst145_p8;
logic [31:0] inst145_p9;
logic [31:0] inst145_p10;
logic [31:0] inst145_p11;
logic [31:0] inst145_p12;
logic [31:0] inst145_p13;
logic [31:0] inst145_p14;
logic [31:0] inst145_p15;
logic [31:0] inst145_p16;
logic [31:0] inst145_p17;
logic [31:0] inst145_p18;
logic [31:0] inst145_p19;
logic [31:0] inst145_p20;
logic [31:0] inst145_p21;
logic [31:0] inst145_p22;
logic [31:0] inst145_p23;
logic [31:0] inst145_p24;
logic [31:0] inst145_p25;
logic [31:0] inst145_p26;
logic [31:0] inst145_p27;
logic [31:0] inst145_p28;
logic [31:0] inst145_p29;
logic [31:0] inst145_p30;
logic [31:0] inst145_p31;
logic [31:0] inst145_p32;
logic [31:0] inst145_p33;
logic [31:0] inst145_p34;
logic [31:0] inst145_p35;
logic [31:0] inst145_p36;
logic [1023:0] inst145_p37;
logic inst145_clk;
logic inst145_reset;
logic [1023:0] inst146_p4;
logic [31:0] inst146_p5;
logic [31:0] inst146_p6;
logic [31:0] inst146_p7;
logic [31:0] inst146_p8;
logic [31:0] inst146_p9;
logic [31:0] inst146_p10;
logic [31:0] inst146_p11;
logic [31:0] inst146_p12;
logic [31:0] inst146_p13;
logic [31:0] inst146_p14;
logic [31:0] inst146_p15;
logic [31:0] inst146_p16;
logic [31:0] inst146_p17;
logic [31:0] inst146_p18;
logic [31:0] inst146_p19;
logic [31:0] inst146_p20;
logic [31:0] inst146_p21;
logic [31:0] inst146_p22;
logic [31:0] inst146_p23;
logic [31:0] inst146_p24;
logic [31:0] inst146_p25;
logic [31:0] inst146_p26;
logic [31:0] inst146_p27;
logic [31:0] inst146_p28;
logic [31:0] inst146_p29;
logic [31:0] inst146_p30;
logic [31:0] inst146_p31;
logic [31:0] inst146_p32;
logic [31:0] inst146_p33;
logic [31:0] inst146_p34;
logic [31:0] inst146_p35;
logic [31:0] inst146_p36;
logic inst146_clk;
logic inst146_reset;
logic [31:0] inst147_p5;
logic [31:0] inst147_p6;
logic [31:0] inst147_p7;
logic [31:0] inst147_p8;
logic [31:0] inst147_p9;
logic [31:0] inst147_p10;
logic [31:0] inst147_p11;
logic [31:0] inst147_p12;
logic [31:0] inst147_p13;
logic [31:0] inst147_p14;
logic [31:0] inst147_p15;
logic [31:0] inst147_p16;
logic [31:0] inst147_p17;
logic [31:0] inst147_p18;
logic [31:0] inst147_p19;
logic [31:0] inst147_p20;
logic [31:0] inst147_p21;
logic [31:0] inst147_p22;
logic [31:0] inst147_p23;
logic [31:0] inst147_p24;
logic [31:0] inst147_p25;
logic [31:0] inst147_p26;
logic [31:0] inst147_p27;
logic [31:0] inst147_p28;
logic [31:0] inst147_p29;
logic [31:0] inst147_p30;
logic [31:0] inst147_p31;
logic [31:0] inst147_p32;
logic [31:0] inst147_p33;
logic [31:0] inst147_p34;
logic [31:0] inst147_p35;
logic [31:0] inst147_p36;
logic [1023:0] inst147_p37;
logic inst147_clk;
logic inst147_reset;
logic [1023:0] inst148_p4;
logic [31:0] inst148_p5;
logic [31:0] inst148_p6;
logic [31:0] inst148_p7;
logic [31:0] inst148_p8;
logic [31:0] inst148_p9;
logic [31:0] inst148_p10;
logic [31:0] inst148_p11;
logic [31:0] inst148_p12;
logic [31:0] inst148_p13;
logic [31:0] inst148_p14;
logic [31:0] inst148_p15;
logic [31:0] inst148_p16;
logic [31:0] inst148_p17;
logic [31:0] inst148_p18;
logic [31:0] inst148_p19;
logic [31:0] inst148_p20;
logic [31:0] inst148_p21;
logic [31:0] inst148_p22;
logic [31:0] inst148_p23;
logic [31:0] inst148_p24;
logic [31:0] inst148_p25;
logic [31:0] inst148_p26;
logic [31:0] inst148_p27;
logic [31:0] inst148_p28;
logic [31:0] inst148_p29;
logic [31:0] inst148_p30;
logic [31:0] inst148_p31;
logic [31:0] inst148_p32;
logic [31:0] inst148_p33;
logic [31:0] inst148_p34;
logic [31:0] inst148_p35;
logic [31:0] inst148_p36;
logic inst148_clk;
logic inst148_reset;
logic [31:0] inst149_p5;
logic [31:0] inst149_p6;
logic [31:0] inst149_p7;
logic [31:0] inst149_p8;
logic [31:0] inst149_p9;
logic [31:0] inst149_p10;
logic [31:0] inst149_p11;
logic [31:0] inst149_p12;
logic [31:0] inst149_p13;
logic [31:0] inst149_p14;
logic [31:0] inst149_p15;
logic [31:0] inst149_p16;
logic [31:0] inst149_p17;
logic [31:0] inst149_p18;
logic [31:0] inst149_p19;
logic [31:0] inst149_p20;
logic [31:0] inst149_p21;
logic [31:0] inst149_p22;
logic [31:0] inst149_p23;
logic [31:0] inst149_p24;
logic [31:0] inst149_p25;
logic [31:0] inst149_p26;
logic [31:0] inst149_p27;
logic [31:0] inst149_p28;
logic [31:0] inst149_p29;
logic [31:0] inst149_p30;
logic [31:0] inst149_p31;
logic [31:0] inst149_p32;
logic [31:0] inst149_p33;
logic [31:0] inst149_p34;
logic [31:0] inst149_p35;
logic [31:0] inst149_p36;
logic [1023:0] inst149_p37;
logic inst149_clk;
logic inst149_reset;
logic [1023:0] inst150_p4;
logic [31:0] inst150_p5;
logic [31:0] inst150_p6;
logic [31:0] inst150_p7;
logic [31:0] inst150_p8;
logic [31:0] inst150_p9;
logic [31:0] inst150_p10;
logic [31:0] inst150_p11;
logic [31:0] inst150_p12;
logic [31:0] inst150_p13;
logic [31:0] inst150_p14;
logic [31:0] inst150_p15;
logic [31:0] inst150_p16;
logic [31:0] inst150_p17;
logic [31:0] inst150_p18;
logic [31:0] inst150_p19;
logic [31:0] inst150_p20;
logic [31:0] inst150_p21;
logic [31:0] inst150_p22;
logic [31:0] inst150_p23;
logic [31:0] inst150_p24;
logic [31:0] inst150_p25;
logic [31:0] inst150_p26;
logic [31:0] inst150_p27;
logic [31:0] inst150_p28;
logic [31:0] inst150_p29;
logic [31:0] inst150_p30;
logic [31:0] inst150_p31;
logic [31:0] inst150_p32;
logic [31:0] inst150_p33;
logic [31:0] inst150_p34;
logic [31:0] inst150_p35;
logic [31:0] inst150_p36;
logic inst150_clk;
logic inst150_reset;
logic [31:0] inst151_p5;
logic [31:0] inst151_p6;
logic [31:0] inst151_p7;
logic [31:0] inst151_p8;
logic [31:0] inst151_p9;
logic [31:0] inst151_p10;
logic [31:0] inst151_p11;
logic [31:0] inst151_p12;
logic [31:0] inst151_p13;
logic [31:0] inst151_p14;
logic [31:0] inst151_p15;
logic [31:0] inst151_p16;
logic [31:0] inst151_p17;
logic [31:0] inst151_p18;
logic [31:0] inst151_p19;
logic [31:0] inst151_p20;
logic [31:0] inst151_p21;
logic [31:0] inst151_p22;
logic [31:0] inst151_p23;
logic [31:0] inst151_p24;
logic [31:0] inst151_p25;
logic [31:0] inst151_p26;
logic [31:0] inst151_p27;
logic [31:0] inst151_p28;
logic [31:0] inst151_p29;
logic [31:0] inst151_p30;
logic [31:0] inst151_p31;
logic [31:0] inst151_p32;
logic [31:0] inst151_p33;
logic [31:0] inst151_p34;
logic [31:0] inst151_p35;
logic [31:0] inst151_p36;
logic [1023:0] inst151_p37;
logic inst151_clk;
logic inst151_reset;
logic [1023:0] inst152_p4;
logic [31:0] inst152_p5;
logic [31:0] inst152_p6;
logic [31:0] inst152_p7;
logic [31:0] inst152_p8;
logic [31:0] inst152_p9;
logic [31:0] inst152_p10;
logic [31:0] inst152_p11;
logic [31:0] inst152_p12;
logic [31:0] inst152_p13;
logic [31:0] inst152_p14;
logic [31:0] inst152_p15;
logic [31:0] inst152_p16;
logic [31:0] inst152_p17;
logic [31:0] inst152_p18;
logic [31:0] inst152_p19;
logic [31:0] inst152_p20;
logic [31:0] inst152_p21;
logic [31:0] inst152_p22;
logic [31:0] inst152_p23;
logic [31:0] inst152_p24;
logic [31:0] inst152_p25;
logic [31:0] inst152_p26;
logic [31:0] inst152_p27;
logic [31:0] inst152_p28;
logic [31:0] inst152_p29;
logic [31:0] inst152_p30;
logic [31:0] inst152_p31;
logic [31:0] inst152_p32;
logic [31:0] inst152_p33;
logic [31:0] inst152_p34;
logic [31:0] inst152_p35;
logic [31:0] inst152_p36;
logic inst152_clk;
logic inst152_reset;
counter_chain_2_52 ev00 (
    ._0_0(ev00__0_0),
    ._0state(ev00__0state),
    ._1_0(ev00__1_0),
    ._1state(ev00__1state),
    .clk(ev00_clk),
    .done(ev00_done),
    .go(ev00_go),
    .reset(ev00_reset)
);
comp35 inst0 (
    .clk(inst0_clk),
    .ev0(inst0_ev0),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
comp48 inst1 (
    .clk(inst1_clk),
    .p17(inst1_p17),
    .p18(inst1_p18),
    .p19(inst1_p19),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .p30(inst1_p30),
    .p31(inst1_p31),
    .p32(inst1_p32),
    .reset(inst1_reset)
);
comp49 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p2(inst2_p2),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p3(inst2_p3),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p38(inst2_p38),
    .p39(inst2_p39),
    .p4(inst2_p4),
    .p40(inst2_p40),
    .p41(inst2_p41),
    .p42(inst2_p42),
    .p43(inst2_p43),
    .p44(inst2_p44),
    .p45(inst2_p45),
    .p46(inst2_p46),
    .p47(inst2_p47),
    .p48(inst2_p48),
    .p49(inst2_p49),
    .p5(inst2_p5),
    .p50(inst2_p50),
    .p51(inst2_p51),
    .p52(inst2_p52),
    .p53(inst2_p53),
    .p54(inst2_p54),
    .p55(inst2_p55),
    .p56(inst2_p56),
    .p57(inst2_p57),
    .p58(inst2_p58),
    .p59(inst2_p59),
    .p6(inst2_p6),
    .p60(inst2_p60),
    .p61(inst2_p61),
    .p62(inst2_p62),
    .p63(inst2_p63),
    .p64(inst2_p64),
    .p65(inst2_p65),
    .p7(inst2_p7),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
comp50 inst3 (
    .clk(inst3_clk),
    .p10(inst3_p10),
    .p11(inst3_p11),
    .p12(inst3_p12),
    .p13(inst3_p13),
    .p14(inst3_p14),
    .p15(inst3_p15),
    .p16(inst3_p16),
    .p17(inst3_p17),
    .p18(inst3_p18),
    .p19(inst3_p19),
    .p2(inst3_p2),
    .p20(inst3_p20),
    .p21(inst3_p21),
    .p22(inst3_p22),
    .p23(inst3_p23),
    .p24(inst3_p24),
    .p25(inst3_p25),
    .p26(inst3_p26),
    .p27(inst3_p27),
    .p28(inst3_p28),
    .p29(inst3_p29),
    .p3(inst3_p3),
    .p30(inst3_p30),
    .p31(inst3_p31),
    .p32(inst3_p32),
    .p33(inst3_p33),
    .p34(inst3_p34),
    .p35(inst3_p35),
    .p36(inst3_p36),
    .p37(inst3_p37),
    .p38(inst3_p38),
    .p39(inst3_p39),
    .p4(inst3_p4),
    .p40(inst3_p40),
    .p41(inst3_p41),
    .p42(inst3_p42),
    .p43(inst3_p43),
    .p44(inst3_p44),
    .p45(inst3_p45),
    .p46(inst3_p46),
    .p47(inst3_p47),
    .p48(inst3_p48),
    .p49(inst3_p49),
    .p5(inst3_p5),
    .p50(inst3_p50),
    .p51(inst3_p51),
    .p52(inst3_p52),
    .p53(inst3_p53),
    .p54(inst3_p54),
    .p55(inst3_p55),
    .p56(inst3_p56),
    .p57(inst3_p57),
    .p58(inst3_p58),
    .p59(inst3_p59),
    .p6(inst3_p6),
    .p60(inst3_p60),
    .p61(inst3_p61),
    .p62(inst3_p62),
    .p63(inst3_p63),
    .p64(inst3_p64),
    .p65(inst3_p65),
    .p7(inst3_p7),
    .p8(inst3_p8),
    .p9(inst3_p9),
    .reset(inst3_reset)
);
Delay # (
    .WIDTH(1024)
) inst4 (
    .clk(inst4_clk),
    .in(inst4_in),
    .out(inst4_out),
    .reset(inst4_reset)
);
comp52 inst5 (
    .clk(inst5_clk),
    .p10(inst5_p10),
    .p11(inst5_p11),
    .p12(inst5_p12),
    .p13(inst5_p13),
    .p14(inst5_p14),
    .p15(inst5_p15),
    .p16(inst5_p16),
    .p17(inst5_p17),
    .p18(inst5_p18),
    .p19(inst5_p19),
    .p2(inst5_p2),
    .p20(inst5_p20),
    .p21(inst5_p21),
    .p22(inst5_p22),
    .p23(inst5_p23),
    .p24(inst5_p24),
    .p25(inst5_p25),
    .p26(inst5_p26),
    .p27(inst5_p27),
    .p28(inst5_p28),
    .p29(inst5_p29),
    .p3(inst5_p3),
    .p30(inst5_p30),
    .p31(inst5_p31),
    .p32(inst5_p32),
    .p33(inst5_p33),
    .p4(inst5_p4),
    .p5(inst5_p5),
    .p6(inst5_p6),
    .p7(inst5_p7),
    .p8(inst5_p8),
    .p9(inst5_p9),
    .reset(inst5_reset)
);
comp53 inst6 (
    .clk(inst6_clk),
    .p10(inst6_p10),
    .p11(inst6_p11),
    .p12(inst6_p12),
    .p13(inst6_p13),
    .p14(inst6_p14),
    .p15(inst6_p15),
    .p16(inst6_p16),
    .p17(inst6_p17),
    .p18(inst6_p18),
    .p19(inst6_p19),
    .p2(inst6_p2),
    .p20(inst6_p20),
    .p21(inst6_p21),
    .p22(inst6_p22),
    .p23(inst6_p23),
    .p24(inst6_p24),
    .p25(inst6_p25),
    .p26(inst6_p26),
    .p27(inst6_p27),
    .p28(inst6_p28),
    .p29(inst6_p29),
    .p3(inst6_p3),
    .p30(inst6_p30),
    .p31(inst6_p31),
    .p32(inst6_p32),
    .p33(inst6_p33),
    .p4(inst6_p4),
    .p5(inst6_p5),
    .p6(inst6_p6),
    .p7(inst6_p7),
    .p8(inst6_p8),
    .p9(inst6_p9),
    .reset(inst6_reset)
);
comp54 inst7 (
    .clk(inst7_clk),
    .p10(inst7_p10),
    .p11(inst7_p11),
    .p12(inst7_p12),
    .p13(inst7_p13),
    .p14(inst7_p14),
    .p15(inst7_p15),
    .p16(inst7_p16),
    .p17(inst7_p17),
    .p18(inst7_p18),
    .p19(inst7_p19),
    .p2(inst7_p2),
    .p20(inst7_p20),
    .p21(inst7_p21),
    .p22(inst7_p22),
    .p23(inst7_p23),
    .p24(inst7_p24),
    .p25(inst7_p25),
    .p26(inst7_p26),
    .p27(inst7_p27),
    .p28(inst7_p28),
    .p29(inst7_p29),
    .p3(inst7_p3),
    .p30(inst7_p30),
    .p31(inst7_p31),
    .p32(inst7_p32),
    .p33(inst7_p33),
    .p4(inst7_p4),
    .p5(inst7_p5),
    .p6(inst7_p6),
    .p7(inst7_p7),
    .p8(inst7_p8),
    .p9(inst7_p9),
    .reset(inst7_reset)
);
comp55 inst8 (
    .clk(inst8_clk),
    .p10(inst8_p10),
    .p11(inst8_p11),
    .p12(inst8_p12),
    .p13(inst8_p13),
    .p14(inst8_p14),
    .p15(inst8_p15),
    .p16(inst8_p16),
    .p17(inst8_p17),
    .p18(inst8_p18),
    .p19(inst8_p19),
    .p2(inst8_p2),
    .p20(inst8_p20),
    .p21(inst8_p21),
    .p22(inst8_p22),
    .p23(inst8_p23),
    .p24(inst8_p24),
    .p25(inst8_p25),
    .p26(inst8_p26),
    .p27(inst8_p27),
    .p28(inst8_p28),
    .p29(inst8_p29),
    .p3(inst8_p3),
    .p30(inst8_p30),
    .p31(inst8_p31),
    .p32(inst8_p32),
    .p33(inst8_p33),
    .p4(inst8_p4),
    .p5(inst8_p5),
    .p6(inst8_p6),
    .p7(inst8_p7),
    .p8(inst8_p8),
    .p9(inst8_p9),
    .reset(inst8_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst9 (
    .clk(inst9_clk),
    .in(inst9_in),
    .out(inst9_out),
    .reset(inst9_reset),
    .write_en(inst9_write_en)
);
comp57 inst10 (
    .clk(inst10_clk),
    .p4(inst10_p4),
    .p5(inst10_p5),
    .p6(inst10_p6),
    .p7(inst10_p7),
    .p8(inst10_p8),
    .reset(inst10_reset)
);
comp63 inst11 (
    .clk(inst11_clk),
    .p5(inst11_p5),
    .p6(inst11_p6),
    .p7(inst11_p7),
    .p8(inst11_p8),
    .p9(inst11_p9),
    .reset(inst11_reset)
);
comp63 inst12 (
    .clk(inst12_clk),
    .p5(inst12_p5),
    .p6(inst12_p6),
    .p7(inst12_p7),
    .p8(inst12_p8),
    .p9(inst12_p9),
    .reset(inst12_reset)
);
comp57 inst13 (
    .clk(inst13_clk),
    .p4(inst13_p4),
    .p5(inst13_p5),
    .p6(inst13_p6),
    .p7(inst13_p7),
    .p8(inst13_p8),
    .reset(inst13_reset)
);
comp57 inst14 (
    .clk(inst14_clk),
    .p4(inst14_p4),
    .p5(inst14_p5),
    .p6(inst14_p6),
    .p7(inst14_p7),
    .p8(inst14_p8),
    .reset(inst14_reset)
);
comp63 inst15 (
    .clk(inst15_clk),
    .p5(inst15_p5),
    .p6(inst15_p6),
    .p7(inst15_p7),
    .p8(inst15_p8),
    .p9(inst15_p9),
    .reset(inst15_reset)
);
comp63 inst16 (
    .clk(inst16_clk),
    .p5(inst16_p5),
    .p6(inst16_p6),
    .p7(inst16_p7),
    .p8(inst16_p8),
    .p9(inst16_p9),
    .reset(inst16_reset)
);
comp57 inst17 (
    .clk(inst17_clk),
    .p4(inst17_p4),
    .p5(inst17_p5),
    .p6(inst17_p6),
    .p7(inst17_p7),
    .p8(inst17_p8),
    .reset(inst17_reset)
);
comp57 inst18 (
    .clk(inst18_clk),
    .p4(inst18_p4),
    .p5(inst18_p5),
    .p6(inst18_p6),
    .p7(inst18_p7),
    .p8(inst18_p8),
    .reset(inst18_reset)
);
comp63 inst19 (
    .clk(inst19_clk),
    .p5(inst19_p5),
    .p6(inst19_p6),
    .p7(inst19_p7),
    .p8(inst19_p8),
    .p9(inst19_p9),
    .reset(inst19_reset)
);
comp63 inst20 (
    .clk(inst20_clk),
    .p5(inst20_p5),
    .p6(inst20_p6),
    .p7(inst20_p7),
    .p8(inst20_p8),
    .p9(inst20_p9),
    .reset(inst20_reset)
);
comp57 inst21 (
    .clk(inst21_clk),
    .p4(inst21_p4),
    .p5(inst21_p5),
    .p6(inst21_p6),
    .p7(inst21_p7),
    .p8(inst21_p8),
    .reset(inst21_reset)
);
comp57 inst22 (
    .clk(inst22_clk),
    .p4(inst22_p4),
    .p5(inst22_p5),
    .p6(inst22_p6),
    .p7(inst22_p7),
    .p8(inst22_p8),
    .reset(inst22_reset)
);
comp63 inst23 (
    .clk(inst23_clk),
    .p5(inst23_p5),
    .p6(inst23_p6),
    .p7(inst23_p7),
    .p8(inst23_p8),
    .p9(inst23_p9),
    .reset(inst23_reset)
);
comp63 inst24 (
    .clk(inst24_clk),
    .p5(inst24_p5),
    .p6(inst24_p6),
    .p7(inst24_p7),
    .p8(inst24_p8),
    .p9(inst24_p9),
    .reset(inst24_reset)
);
comp57 inst25 (
    .clk(inst25_clk),
    .p4(inst25_p4),
    .p5(inst25_p5),
    .p6(inst25_p6),
    .p7(inst25_p7),
    .p8(inst25_p8),
    .reset(inst25_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst26 (
    .clk(inst26_clk),
    .in(inst26_in),
    .out(inst26_out),
    .reset(inst26_reset),
    .write_en(inst26_write_en)
);
comp57 inst27 (
    .clk(inst27_clk),
    .p4(inst27_p4),
    .p5(inst27_p5),
    .p6(inst27_p6),
    .p7(inst27_p7),
    .p8(inst27_p8),
    .reset(inst27_reset)
);
comp63 inst28 (
    .clk(inst28_clk),
    .p5(inst28_p5),
    .p6(inst28_p6),
    .p7(inst28_p7),
    .p8(inst28_p8),
    .p9(inst28_p9),
    .reset(inst28_reset)
);
comp63 inst29 (
    .clk(inst29_clk),
    .p5(inst29_p5),
    .p6(inst29_p6),
    .p7(inst29_p7),
    .p8(inst29_p8),
    .p9(inst29_p9),
    .reset(inst29_reset)
);
comp57 inst30 (
    .clk(inst30_clk),
    .p4(inst30_p4),
    .p5(inst30_p5),
    .p6(inst30_p6),
    .p7(inst30_p7),
    .p8(inst30_p8),
    .reset(inst30_reset)
);
comp57 inst31 (
    .clk(inst31_clk),
    .p4(inst31_p4),
    .p5(inst31_p5),
    .p6(inst31_p6),
    .p7(inst31_p7),
    .p8(inst31_p8),
    .reset(inst31_reset)
);
comp63 inst32 (
    .clk(inst32_clk),
    .p5(inst32_p5),
    .p6(inst32_p6),
    .p7(inst32_p7),
    .p8(inst32_p8),
    .p9(inst32_p9),
    .reset(inst32_reset)
);
comp63 inst33 (
    .clk(inst33_clk),
    .p5(inst33_p5),
    .p6(inst33_p6),
    .p7(inst33_p7),
    .p8(inst33_p8),
    .p9(inst33_p9),
    .reset(inst33_reset)
);
comp57 inst34 (
    .clk(inst34_clk),
    .p4(inst34_p4),
    .p5(inst34_p5),
    .p6(inst34_p6),
    .p7(inst34_p7),
    .p8(inst34_p8),
    .reset(inst34_reset)
);
comp57 inst35 (
    .clk(inst35_clk),
    .p4(inst35_p4),
    .p5(inst35_p5),
    .p6(inst35_p6),
    .p7(inst35_p7),
    .p8(inst35_p8),
    .reset(inst35_reset)
);
comp63 inst36 (
    .clk(inst36_clk),
    .p5(inst36_p5),
    .p6(inst36_p6),
    .p7(inst36_p7),
    .p8(inst36_p8),
    .p9(inst36_p9),
    .reset(inst36_reset)
);
comp63 inst37 (
    .clk(inst37_clk),
    .p5(inst37_p5),
    .p6(inst37_p6),
    .p7(inst37_p7),
    .p8(inst37_p8),
    .p9(inst37_p9),
    .reset(inst37_reset)
);
comp57 inst38 (
    .clk(inst38_clk),
    .p4(inst38_p4),
    .p5(inst38_p5),
    .p6(inst38_p6),
    .p7(inst38_p7),
    .p8(inst38_p8),
    .reset(inst38_reset)
);
comp57 inst39 (
    .clk(inst39_clk),
    .p4(inst39_p4),
    .p5(inst39_p5),
    .p6(inst39_p6),
    .p7(inst39_p7),
    .p8(inst39_p8),
    .reset(inst39_reset)
);
comp63 inst40 (
    .clk(inst40_clk),
    .p5(inst40_p5),
    .p6(inst40_p6),
    .p7(inst40_p7),
    .p8(inst40_p8),
    .p9(inst40_p9),
    .reset(inst40_reset)
);
comp63 inst41 (
    .clk(inst41_clk),
    .p5(inst41_p5),
    .p6(inst41_p6),
    .p7(inst41_p7),
    .p8(inst41_p8),
    .p9(inst41_p9),
    .reset(inst41_reset)
);
comp57 inst42 (
    .clk(inst42_clk),
    .p4(inst42_p4),
    .p5(inst42_p5),
    .p6(inst42_p6),
    .p7(inst42_p7),
    .p8(inst42_p8),
    .reset(inst42_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst43 (
    .clk(inst43_clk),
    .in(inst43_in),
    .out(inst43_out),
    .reset(inst43_reset),
    .write_en(inst43_write_en)
);
comp57 inst44 (
    .clk(inst44_clk),
    .p4(inst44_p4),
    .p5(inst44_p5),
    .p6(inst44_p6),
    .p7(inst44_p7),
    .p8(inst44_p8),
    .reset(inst44_reset)
);
comp63 inst45 (
    .clk(inst45_clk),
    .p5(inst45_p5),
    .p6(inst45_p6),
    .p7(inst45_p7),
    .p8(inst45_p8),
    .p9(inst45_p9),
    .reset(inst45_reset)
);
comp63 inst46 (
    .clk(inst46_clk),
    .p5(inst46_p5),
    .p6(inst46_p6),
    .p7(inst46_p7),
    .p8(inst46_p8),
    .p9(inst46_p9),
    .reset(inst46_reset)
);
comp57 inst47 (
    .clk(inst47_clk),
    .p4(inst47_p4),
    .p5(inst47_p5),
    .p6(inst47_p6),
    .p7(inst47_p7),
    .p8(inst47_p8),
    .reset(inst47_reset)
);
comp57 inst48 (
    .clk(inst48_clk),
    .p4(inst48_p4),
    .p5(inst48_p5),
    .p6(inst48_p6),
    .p7(inst48_p7),
    .p8(inst48_p8),
    .reset(inst48_reset)
);
comp63 inst49 (
    .clk(inst49_clk),
    .p5(inst49_p5),
    .p6(inst49_p6),
    .p7(inst49_p7),
    .p8(inst49_p8),
    .p9(inst49_p9),
    .reset(inst49_reset)
);
comp63 inst50 (
    .clk(inst50_clk),
    .p5(inst50_p5),
    .p6(inst50_p6),
    .p7(inst50_p7),
    .p8(inst50_p8),
    .p9(inst50_p9),
    .reset(inst50_reset)
);
comp57 inst51 (
    .clk(inst51_clk),
    .p4(inst51_p4),
    .p5(inst51_p5),
    .p6(inst51_p6),
    .p7(inst51_p7),
    .p8(inst51_p8),
    .reset(inst51_reset)
);
comp57 inst52 (
    .clk(inst52_clk),
    .p4(inst52_p4),
    .p5(inst52_p5),
    .p6(inst52_p6),
    .p7(inst52_p7),
    .p8(inst52_p8),
    .reset(inst52_reset)
);
comp63 inst53 (
    .clk(inst53_clk),
    .p5(inst53_p5),
    .p6(inst53_p6),
    .p7(inst53_p7),
    .p8(inst53_p8),
    .p9(inst53_p9),
    .reset(inst53_reset)
);
comp63 inst54 (
    .clk(inst54_clk),
    .p5(inst54_p5),
    .p6(inst54_p6),
    .p7(inst54_p7),
    .p8(inst54_p8),
    .p9(inst54_p9),
    .reset(inst54_reset)
);
comp57 inst55 (
    .clk(inst55_clk),
    .p4(inst55_p4),
    .p5(inst55_p5),
    .p6(inst55_p6),
    .p7(inst55_p7),
    .p8(inst55_p8),
    .reset(inst55_reset)
);
comp57 inst56 (
    .clk(inst56_clk),
    .p4(inst56_p4),
    .p5(inst56_p5),
    .p6(inst56_p6),
    .p7(inst56_p7),
    .p8(inst56_p8),
    .reset(inst56_reset)
);
comp63 inst57 (
    .clk(inst57_clk),
    .p5(inst57_p5),
    .p6(inst57_p6),
    .p7(inst57_p7),
    .p8(inst57_p8),
    .p9(inst57_p9),
    .reset(inst57_reset)
);
comp63 inst58 (
    .clk(inst58_clk),
    .p5(inst58_p5),
    .p6(inst58_p6),
    .p7(inst58_p7),
    .p8(inst58_p8),
    .p9(inst58_p9),
    .reset(inst58_reset)
);
comp57 inst59 (
    .clk(inst59_clk),
    .p4(inst59_p4),
    .p5(inst59_p5),
    .p6(inst59_p6),
    .p7(inst59_p7),
    .p8(inst59_p8),
    .reset(inst59_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst60 (
    .clk(inst60_clk),
    .in(inst60_in),
    .out(inst60_out),
    .reset(inst60_reset),
    .write_en(inst60_write_en)
);
comp57 inst61 (
    .clk(inst61_clk),
    .p4(inst61_p4),
    .p5(inst61_p5),
    .p6(inst61_p6),
    .p7(inst61_p7),
    .p8(inst61_p8),
    .reset(inst61_reset)
);
comp63 inst62 (
    .clk(inst62_clk),
    .p5(inst62_p5),
    .p6(inst62_p6),
    .p7(inst62_p7),
    .p8(inst62_p8),
    .p9(inst62_p9),
    .reset(inst62_reset)
);
comp63 inst63 (
    .clk(inst63_clk),
    .p5(inst63_p5),
    .p6(inst63_p6),
    .p7(inst63_p7),
    .p8(inst63_p8),
    .p9(inst63_p9),
    .reset(inst63_reset)
);
comp57 inst64 (
    .clk(inst64_clk),
    .p4(inst64_p4),
    .p5(inst64_p5),
    .p6(inst64_p6),
    .p7(inst64_p7),
    .p8(inst64_p8),
    .reset(inst64_reset)
);
comp57 inst65 (
    .clk(inst65_clk),
    .p4(inst65_p4),
    .p5(inst65_p5),
    .p6(inst65_p6),
    .p7(inst65_p7),
    .p8(inst65_p8),
    .reset(inst65_reset)
);
comp63 inst66 (
    .clk(inst66_clk),
    .p5(inst66_p5),
    .p6(inst66_p6),
    .p7(inst66_p7),
    .p8(inst66_p8),
    .p9(inst66_p9),
    .reset(inst66_reset)
);
comp63 inst67 (
    .clk(inst67_clk),
    .p5(inst67_p5),
    .p6(inst67_p6),
    .p7(inst67_p7),
    .p8(inst67_p8),
    .p9(inst67_p9),
    .reset(inst67_reset)
);
comp57 inst68 (
    .clk(inst68_clk),
    .p4(inst68_p4),
    .p5(inst68_p5),
    .p6(inst68_p6),
    .p7(inst68_p7),
    .p8(inst68_p8),
    .reset(inst68_reset)
);
comp57 inst69 (
    .clk(inst69_clk),
    .p4(inst69_p4),
    .p5(inst69_p5),
    .p6(inst69_p6),
    .p7(inst69_p7),
    .p8(inst69_p8),
    .reset(inst69_reset)
);
comp63 inst70 (
    .clk(inst70_clk),
    .p5(inst70_p5),
    .p6(inst70_p6),
    .p7(inst70_p7),
    .p8(inst70_p8),
    .p9(inst70_p9),
    .reset(inst70_reset)
);
comp63 inst71 (
    .clk(inst71_clk),
    .p5(inst71_p5),
    .p6(inst71_p6),
    .p7(inst71_p7),
    .p8(inst71_p8),
    .p9(inst71_p9),
    .reset(inst71_reset)
);
comp57 inst72 (
    .clk(inst72_clk),
    .p4(inst72_p4),
    .p5(inst72_p5),
    .p6(inst72_p6),
    .p7(inst72_p7),
    .p8(inst72_p8),
    .reset(inst72_reset)
);
comp57 inst73 (
    .clk(inst73_clk),
    .p4(inst73_p4),
    .p5(inst73_p5),
    .p6(inst73_p6),
    .p7(inst73_p7),
    .p8(inst73_p8),
    .reset(inst73_reset)
);
comp63 inst74 (
    .clk(inst74_clk),
    .p5(inst74_p5),
    .p6(inst74_p6),
    .p7(inst74_p7),
    .p8(inst74_p8),
    .p9(inst74_p9),
    .reset(inst74_reset)
);
comp63 inst75 (
    .clk(inst75_clk),
    .p5(inst75_p5),
    .p6(inst75_p6),
    .p7(inst75_p7),
    .p8(inst75_p8),
    .p9(inst75_p9),
    .reset(inst75_reset)
);
comp57 inst76 (
    .clk(inst76_clk),
    .p4(inst76_p4),
    .p5(inst76_p5),
    .p6(inst76_p6),
    .p7(inst76_p7),
    .p8(inst76_p8),
    .reset(inst76_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst77 (
    .clk(inst77_clk),
    .in(inst77_in),
    .out(inst77_out),
    .reset(inst77_reset),
    .write_en(inst77_write_en)
);
comp57 inst78 (
    .clk(inst78_clk),
    .p4(inst78_p4),
    .p5(inst78_p5),
    .p6(inst78_p6),
    .p7(inst78_p7),
    .p8(inst78_p8),
    .reset(inst78_reset)
);
comp63 inst79 (
    .clk(inst79_clk),
    .p5(inst79_p5),
    .p6(inst79_p6),
    .p7(inst79_p7),
    .p8(inst79_p8),
    .p9(inst79_p9),
    .reset(inst79_reset)
);
comp63 inst80 (
    .clk(inst80_clk),
    .p5(inst80_p5),
    .p6(inst80_p6),
    .p7(inst80_p7),
    .p8(inst80_p8),
    .p9(inst80_p9),
    .reset(inst80_reset)
);
comp57 inst81 (
    .clk(inst81_clk),
    .p4(inst81_p4),
    .p5(inst81_p5),
    .p6(inst81_p6),
    .p7(inst81_p7),
    .p8(inst81_p8),
    .reset(inst81_reset)
);
comp57 inst82 (
    .clk(inst82_clk),
    .p4(inst82_p4),
    .p5(inst82_p5),
    .p6(inst82_p6),
    .p7(inst82_p7),
    .p8(inst82_p8),
    .reset(inst82_reset)
);
comp63 inst83 (
    .clk(inst83_clk),
    .p5(inst83_p5),
    .p6(inst83_p6),
    .p7(inst83_p7),
    .p8(inst83_p8),
    .p9(inst83_p9),
    .reset(inst83_reset)
);
comp63 inst84 (
    .clk(inst84_clk),
    .p5(inst84_p5),
    .p6(inst84_p6),
    .p7(inst84_p7),
    .p8(inst84_p8),
    .p9(inst84_p9),
    .reset(inst84_reset)
);
comp57 inst85 (
    .clk(inst85_clk),
    .p4(inst85_p4),
    .p5(inst85_p5),
    .p6(inst85_p6),
    .p7(inst85_p7),
    .p8(inst85_p8),
    .reset(inst85_reset)
);
comp57 inst86 (
    .clk(inst86_clk),
    .p4(inst86_p4),
    .p5(inst86_p5),
    .p6(inst86_p6),
    .p7(inst86_p7),
    .p8(inst86_p8),
    .reset(inst86_reset)
);
comp63 inst87 (
    .clk(inst87_clk),
    .p5(inst87_p5),
    .p6(inst87_p6),
    .p7(inst87_p7),
    .p8(inst87_p8),
    .p9(inst87_p9),
    .reset(inst87_reset)
);
comp63 inst88 (
    .clk(inst88_clk),
    .p5(inst88_p5),
    .p6(inst88_p6),
    .p7(inst88_p7),
    .p8(inst88_p8),
    .p9(inst88_p9),
    .reset(inst88_reset)
);
comp57 inst89 (
    .clk(inst89_clk),
    .p4(inst89_p4),
    .p5(inst89_p5),
    .p6(inst89_p6),
    .p7(inst89_p7),
    .p8(inst89_p8),
    .reset(inst89_reset)
);
comp57 inst90 (
    .clk(inst90_clk),
    .p4(inst90_p4),
    .p5(inst90_p5),
    .p6(inst90_p6),
    .p7(inst90_p7),
    .p8(inst90_p8),
    .reset(inst90_reset)
);
comp63 inst91 (
    .clk(inst91_clk),
    .p5(inst91_p5),
    .p6(inst91_p6),
    .p7(inst91_p7),
    .p8(inst91_p8),
    .p9(inst91_p9),
    .reset(inst91_reset)
);
comp63 inst92 (
    .clk(inst92_clk),
    .p5(inst92_p5),
    .p6(inst92_p6),
    .p7(inst92_p7),
    .p8(inst92_p8),
    .p9(inst92_p9),
    .reset(inst92_reset)
);
comp57 inst93 (
    .clk(inst93_clk),
    .p4(inst93_p4),
    .p5(inst93_p5),
    .p6(inst93_p6),
    .p7(inst93_p7),
    .p8(inst93_p8),
    .reset(inst93_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst94 (
    .clk(inst94_clk),
    .in(inst94_in),
    .out(inst94_out),
    .reset(inst94_reset),
    .write_en(inst94_write_en)
);
comp57 inst95 (
    .clk(inst95_clk),
    .p4(inst95_p4),
    .p5(inst95_p5),
    .p6(inst95_p6),
    .p7(inst95_p7),
    .p8(inst95_p8),
    .reset(inst95_reset)
);
comp63 inst96 (
    .clk(inst96_clk),
    .p5(inst96_p5),
    .p6(inst96_p6),
    .p7(inst96_p7),
    .p8(inst96_p8),
    .p9(inst96_p9),
    .reset(inst96_reset)
);
comp63 inst97 (
    .clk(inst97_clk),
    .p5(inst97_p5),
    .p6(inst97_p6),
    .p7(inst97_p7),
    .p8(inst97_p8),
    .p9(inst97_p9),
    .reset(inst97_reset)
);
comp57 inst98 (
    .clk(inst98_clk),
    .p4(inst98_p4),
    .p5(inst98_p5),
    .p6(inst98_p6),
    .p7(inst98_p7),
    .p8(inst98_p8),
    .reset(inst98_reset)
);
comp57 inst99 (
    .clk(inst99_clk),
    .p4(inst99_p4),
    .p5(inst99_p5),
    .p6(inst99_p6),
    .p7(inst99_p7),
    .p8(inst99_p8),
    .reset(inst99_reset)
);
comp63 inst100 (
    .clk(inst100_clk),
    .p5(inst100_p5),
    .p6(inst100_p6),
    .p7(inst100_p7),
    .p8(inst100_p8),
    .p9(inst100_p9),
    .reset(inst100_reset)
);
comp63 inst101 (
    .clk(inst101_clk),
    .p5(inst101_p5),
    .p6(inst101_p6),
    .p7(inst101_p7),
    .p8(inst101_p8),
    .p9(inst101_p9),
    .reset(inst101_reset)
);
comp57 inst102 (
    .clk(inst102_clk),
    .p4(inst102_p4),
    .p5(inst102_p5),
    .p6(inst102_p6),
    .p7(inst102_p7),
    .p8(inst102_p8),
    .reset(inst102_reset)
);
comp57 inst103 (
    .clk(inst103_clk),
    .p4(inst103_p4),
    .p5(inst103_p5),
    .p6(inst103_p6),
    .p7(inst103_p7),
    .p8(inst103_p8),
    .reset(inst103_reset)
);
comp63 inst104 (
    .clk(inst104_clk),
    .p5(inst104_p5),
    .p6(inst104_p6),
    .p7(inst104_p7),
    .p8(inst104_p8),
    .p9(inst104_p9),
    .reset(inst104_reset)
);
comp63 inst105 (
    .clk(inst105_clk),
    .p5(inst105_p5),
    .p6(inst105_p6),
    .p7(inst105_p7),
    .p8(inst105_p8),
    .p9(inst105_p9),
    .reset(inst105_reset)
);
comp57 inst106 (
    .clk(inst106_clk),
    .p4(inst106_p4),
    .p5(inst106_p5),
    .p6(inst106_p6),
    .p7(inst106_p7),
    .p8(inst106_p8),
    .reset(inst106_reset)
);
comp57 inst107 (
    .clk(inst107_clk),
    .p4(inst107_p4),
    .p5(inst107_p5),
    .p6(inst107_p6),
    .p7(inst107_p7),
    .p8(inst107_p8),
    .reset(inst107_reset)
);
comp63 inst108 (
    .clk(inst108_clk),
    .p5(inst108_p5),
    .p6(inst108_p6),
    .p7(inst108_p7),
    .p8(inst108_p8),
    .p9(inst108_p9),
    .reset(inst108_reset)
);
comp63 inst109 (
    .clk(inst109_clk),
    .p5(inst109_p5),
    .p6(inst109_p6),
    .p7(inst109_p7),
    .p8(inst109_p8),
    .p9(inst109_p9),
    .reset(inst109_reset)
);
comp57 inst110 (
    .clk(inst110_clk),
    .p4(inst110_p4),
    .p5(inst110_p5),
    .p6(inst110_p6),
    .p7(inst110_p7),
    .p8(inst110_p8),
    .reset(inst110_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst111 (
    .clk(inst111_clk),
    .in(inst111_in),
    .out(inst111_out),
    .reset(inst111_reset),
    .write_en(inst111_write_en)
);
comp57 inst112 (
    .clk(inst112_clk),
    .p4(inst112_p4),
    .p5(inst112_p5),
    .p6(inst112_p6),
    .p7(inst112_p7),
    .p8(inst112_p8),
    .reset(inst112_reset)
);
comp63 inst113 (
    .clk(inst113_clk),
    .p5(inst113_p5),
    .p6(inst113_p6),
    .p7(inst113_p7),
    .p8(inst113_p8),
    .p9(inst113_p9),
    .reset(inst113_reset)
);
comp63 inst114 (
    .clk(inst114_clk),
    .p5(inst114_p5),
    .p6(inst114_p6),
    .p7(inst114_p7),
    .p8(inst114_p8),
    .p9(inst114_p9),
    .reset(inst114_reset)
);
comp57 inst115 (
    .clk(inst115_clk),
    .p4(inst115_p4),
    .p5(inst115_p5),
    .p6(inst115_p6),
    .p7(inst115_p7),
    .p8(inst115_p8),
    .reset(inst115_reset)
);
comp57 inst116 (
    .clk(inst116_clk),
    .p4(inst116_p4),
    .p5(inst116_p5),
    .p6(inst116_p6),
    .p7(inst116_p7),
    .p8(inst116_p8),
    .reset(inst116_reset)
);
comp63 inst117 (
    .clk(inst117_clk),
    .p5(inst117_p5),
    .p6(inst117_p6),
    .p7(inst117_p7),
    .p8(inst117_p8),
    .p9(inst117_p9),
    .reset(inst117_reset)
);
comp63 inst118 (
    .clk(inst118_clk),
    .p5(inst118_p5),
    .p6(inst118_p6),
    .p7(inst118_p7),
    .p8(inst118_p8),
    .p9(inst118_p9),
    .reset(inst118_reset)
);
comp57 inst119 (
    .clk(inst119_clk),
    .p4(inst119_p4),
    .p5(inst119_p5),
    .p6(inst119_p6),
    .p7(inst119_p7),
    .p8(inst119_p8),
    .reset(inst119_reset)
);
comp57 inst120 (
    .clk(inst120_clk),
    .p4(inst120_p4),
    .p5(inst120_p5),
    .p6(inst120_p6),
    .p7(inst120_p7),
    .p8(inst120_p8),
    .reset(inst120_reset)
);
comp63 inst121 (
    .clk(inst121_clk),
    .p5(inst121_p5),
    .p6(inst121_p6),
    .p7(inst121_p7),
    .p8(inst121_p8),
    .p9(inst121_p9),
    .reset(inst121_reset)
);
comp63 inst122 (
    .clk(inst122_clk),
    .p5(inst122_p5),
    .p6(inst122_p6),
    .p7(inst122_p7),
    .p8(inst122_p8),
    .p9(inst122_p9),
    .reset(inst122_reset)
);
comp57 inst123 (
    .clk(inst123_clk),
    .p4(inst123_p4),
    .p5(inst123_p5),
    .p6(inst123_p6),
    .p7(inst123_p7),
    .p8(inst123_p8),
    .reset(inst123_reset)
);
comp57 inst124 (
    .clk(inst124_clk),
    .p4(inst124_p4),
    .p5(inst124_p5),
    .p6(inst124_p6),
    .p7(inst124_p7),
    .p8(inst124_p8),
    .reset(inst124_reset)
);
comp63 inst125 (
    .clk(inst125_clk),
    .p5(inst125_p5),
    .p6(inst125_p6),
    .p7(inst125_p7),
    .p8(inst125_p8),
    .p9(inst125_p9),
    .reset(inst125_reset)
);
comp63 inst126 (
    .clk(inst126_clk),
    .p5(inst126_p5),
    .p6(inst126_p6),
    .p7(inst126_p7),
    .p8(inst126_p8),
    .p9(inst126_p9),
    .reset(inst126_reset)
);
comp57 inst127 (
    .clk(inst127_clk),
    .p4(inst127_p4),
    .p5(inst127_p5),
    .p6(inst127_p6),
    .p7(inst127_p7),
    .p8(inst127_p8),
    .reset(inst127_reset)
);
PassThroughRegister # (
    .WIDTH(128)
) inst128 (
    .clk(inst128_clk),
    .in(inst128_in),
    .out(inst128_out),
    .reset(inst128_reset),
    .write_en(inst128_write_en)
);
comp57 inst129 (
    .clk(inst129_clk),
    .p4(inst129_p4),
    .p5(inst129_p5),
    .p6(inst129_p6),
    .p7(inst129_p7),
    .p8(inst129_p8),
    .reset(inst129_reset)
);
comp63 inst130 (
    .clk(inst130_clk),
    .p5(inst130_p5),
    .p6(inst130_p6),
    .p7(inst130_p7),
    .p8(inst130_p8),
    .p9(inst130_p9),
    .reset(inst130_reset)
);
comp63 inst131 (
    .clk(inst131_clk),
    .p5(inst131_p5),
    .p6(inst131_p6),
    .p7(inst131_p7),
    .p8(inst131_p8),
    .p9(inst131_p9),
    .reset(inst131_reset)
);
comp57 inst132 (
    .clk(inst132_clk),
    .p4(inst132_p4),
    .p5(inst132_p5),
    .p6(inst132_p6),
    .p7(inst132_p7),
    .p8(inst132_p8),
    .reset(inst132_reset)
);
comp57 inst133 (
    .clk(inst133_clk),
    .p4(inst133_p4),
    .p5(inst133_p5),
    .p6(inst133_p6),
    .p7(inst133_p7),
    .p8(inst133_p8),
    .reset(inst133_reset)
);
comp63 inst134 (
    .clk(inst134_clk),
    .p5(inst134_p5),
    .p6(inst134_p6),
    .p7(inst134_p7),
    .p8(inst134_p8),
    .p9(inst134_p9),
    .reset(inst134_reset)
);
comp63 inst135 (
    .clk(inst135_clk),
    .p5(inst135_p5),
    .p6(inst135_p6),
    .p7(inst135_p7),
    .p8(inst135_p8),
    .p9(inst135_p9),
    .reset(inst135_reset)
);
comp57 inst136 (
    .clk(inst136_clk),
    .p4(inst136_p4),
    .p5(inst136_p5),
    .p6(inst136_p6),
    .p7(inst136_p7),
    .p8(inst136_p8),
    .reset(inst136_reset)
);
comp57 inst137 (
    .clk(inst137_clk),
    .p4(inst137_p4),
    .p5(inst137_p5),
    .p6(inst137_p6),
    .p7(inst137_p7),
    .p8(inst137_p8),
    .reset(inst137_reset)
);
comp63 inst138 (
    .clk(inst138_clk),
    .p5(inst138_p5),
    .p6(inst138_p6),
    .p7(inst138_p7),
    .p8(inst138_p8),
    .p9(inst138_p9),
    .reset(inst138_reset)
);
comp63 inst139 (
    .clk(inst139_clk),
    .p5(inst139_p5),
    .p6(inst139_p6),
    .p7(inst139_p7),
    .p8(inst139_p8),
    .p9(inst139_p9),
    .reset(inst139_reset)
);
comp57 inst140 (
    .clk(inst140_clk),
    .p4(inst140_p4),
    .p5(inst140_p5),
    .p6(inst140_p6),
    .p7(inst140_p7),
    .p8(inst140_p8),
    .reset(inst140_reset)
);
comp57 inst141 (
    .clk(inst141_clk),
    .p4(inst141_p4),
    .p5(inst141_p5),
    .p6(inst141_p6),
    .p7(inst141_p7),
    .p8(inst141_p8),
    .reset(inst141_reset)
);
comp63 inst142 (
    .clk(inst142_clk),
    .p5(inst142_p5),
    .p6(inst142_p6),
    .p7(inst142_p7),
    .p8(inst142_p8),
    .p9(inst142_p9),
    .reset(inst142_reset)
);
comp63 inst143 (
    .clk(inst143_clk),
    .p5(inst143_p5),
    .p6(inst143_p6),
    .p7(inst143_p7),
    .p8(inst143_p8),
    .p9(inst143_p9),
    .reset(inst143_reset)
);
comp57 inst144 (
    .clk(inst144_clk),
    .p4(inst144_p4),
    .p5(inst144_p5),
    .p6(inst144_p6),
    .p7(inst144_p7),
    .p8(inst144_p8),
    .reset(inst144_reset)
);
comp92 inst145 (
    .clk(inst145_clk),
    .p10(inst145_p10),
    .p11(inst145_p11),
    .p12(inst145_p12),
    .p13(inst145_p13),
    .p14(inst145_p14),
    .p15(inst145_p15),
    .p16(inst145_p16),
    .p17(inst145_p17),
    .p18(inst145_p18),
    .p19(inst145_p19),
    .p20(inst145_p20),
    .p21(inst145_p21),
    .p22(inst145_p22),
    .p23(inst145_p23),
    .p24(inst145_p24),
    .p25(inst145_p25),
    .p26(inst145_p26),
    .p27(inst145_p27),
    .p28(inst145_p28),
    .p29(inst145_p29),
    .p30(inst145_p30),
    .p31(inst145_p31),
    .p32(inst145_p32),
    .p33(inst145_p33),
    .p34(inst145_p34),
    .p35(inst145_p35),
    .p36(inst145_p36),
    .p37(inst145_p37),
    .p5(inst145_p5),
    .p6(inst145_p6),
    .p7(inst145_p7),
    .p8(inst145_p8),
    .p9(inst145_p9),
    .reset(inst145_reset)
);
comp93 inst146 (
    .clk(inst146_clk),
    .p10(inst146_p10),
    .p11(inst146_p11),
    .p12(inst146_p12),
    .p13(inst146_p13),
    .p14(inst146_p14),
    .p15(inst146_p15),
    .p16(inst146_p16),
    .p17(inst146_p17),
    .p18(inst146_p18),
    .p19(inst146_p19),
    .p20(inst146_p20),
    .p21(inst146_p21),
    .p22(inst146_p22),
    .p23(inst146_p23),
    .p24(inst146_p24),
    .p25(inst146_p25),
    .p26(inst146_p26),
    .p27(inst146_p27),
    .p28(inst146_p28),
    .p29(inst146_p29),
    .p30(inst146_p30),
    .p31(inst146_p31),
    .p32(inst146_p32),
    .p33(inst146_p33),
    .p34(inst146_p34),
    .p35(inst146_p35),
    .p36(inst146_p36),
    .p4(inst146_p4),
    .p5(inst146_p5),
    .p6(inst146_p6),
    .p7(inst146_p7),
    .p8(inst146_p8),
    .p9(inst146_p9),
    .reset(inst146_reset)
);
comp92 inst147 (
    .clk(inst147_clk),
    .p10(inst147_p10),
    .p11(inst147_p11),
    .p12(inst147_p12),
    .p13(inst147_p13),
    .p14(inst147_p14),
    .p15(inst147_p15),
    .p16(inst147_p16),
    .p17(inst147_p17),
    .p18(inst147_p18),
    .p19(inst147_p19),
    .p20(inst147_p20),
    .p21(inst147_p21),
    .p22(inst147_p22),
    .p23(inst147_p23),
    .p24(inst147_p24),
    .p25(inst147_p25),
    .p26(inst147_p26),
    .p27(inst147_p27),
    .p28(inst147_p28),
    .p29(inst147_p29),
    .p30(inst147_p30),
    .p31(inst147_p31),
    .p32(inst147_p32),
    .p33(inst147_p33),
    .p34(inst147_p34),
    .p35(inst147_p35),
    .p36(inst147_p36),
    .p37(inst147_p37),
    .p5(inst147_p5),
    .p6(inst147_p6),
    .p7(inst147_p7),
    .p8(inst147_p8),
    .p9(inst147_p9),
    .reset(inst147_reset)
);
comp93 inst148 (
    .clk(inst148_clk),
    .p10(inst148_p10),
    .p11(inst148_p11),
    .p12(inst148_p12),
    .p13(inst148_p13),
    .p14(inst148_p14),
    .p15(inst148_p15),
    .p16(inst148_p16),
    .p17(inst148_p17),
    .p18(inst148_p18),
    .p19(inst148_p19),
    .p20(inst148_p20),
    .p21(inst148_p21),
    .p22(inst148_p22),
    .p23(inst148_p23),
    .p24(inst148_p24),
    .p25(inst148_p25),
    .p26(inst148_p26),
    .p27(inst148_p27),
    .p28(inst148_p28),
    .p29(inst148_p29),
    .p30(inst148_p30),
    .p31(inst148_p31),
    .p32(inst148_p32),
    .p33(inst148_p33),
    .p34(inst148_p34),
    .p35(inst148_p35),
    .p36(inst148_p36),
    .p4(inst148_p4),
    .p5(inst148_p5),
    .p6(inst148_p6),
    .p7(inst148_p7),
    .p8(inst148_p8),
    .p9(inst148_p9),
    .reset(inst148_reset)
);
comp92 inst149 (
    .clk(inst149_clk),
    .p10(inst149_p10),
    .p11(inst149_p11),
    .p12(inst149_p12),
    .p13(inst149_p13),
    .p14(inst149_p14),
    .p15(inst149_p15),
    .p16(inst149_p16),
    .p17(inst149_p17),
    .p18(inst149_p18),
    .p19(inst149_p19),
    .p20(inst149_p20),
    .p21(inst149_p21),
    .p22(inst149_p22),
    .p23(inst149_p23),
    .p24(inst149_p24),
    .p25(inst149_p25),
    .p26(inst149_p26),
    .p27(inst149_p27),
    .p28(inst149_p28),
    .p29(inst149_p29),
    .p30(inst149_p30),
    .p31(inst149_p31),
    .p32(inst149_p32),
    .p33(inst149_p33),
    .p34(inst149_p34),
    .p35(inst149_p35),
    .p36(inst149_p36),
    .p37(inst149_p37),
    .p5(inst149_p5),
    .p6(inst149_p6),
    .p7(inst149_p7),
    .p8(inst149_p8),
    .p9(inst149_p9),
    .reset(inst149_reset)
);
comp93 inst150 (
    .clk(inst150_clk),
    .p10(inst150_p10),
    .p11(inst150_p11),
    .p12(inst150_p12),
    .p13(inst150_p13),
    .p14(inst150_p14),
    .p15(inst150_p15),
    .p16(inst150_p16),
    .p17(inst150_p17),
    .p18(inst150_p18),
    .p19(inst150_p19),
    .p20(inst150_p20),
    .p21(inst150_p21),
    .p22(inst150_p22),
    .p23(inst150_p23),
    .p24(inst150_p24),
    .p25(inst150_p25),
    .p26(inst150_p26),
    .p27(inst150_p27),
    .p28(inst150_p28),
    .p29(inst150_p29),
    .p30(inst150_p30),
    .p31(inst150_p31),
    .p32(inst150_p32),
    .p33(inst150_p33),
    .p34(inst150_p34),
    .p35(inst150_p35),
    .p36(inst150_p36),
    .p4(inst150_p4),
    .p5(inst150_p5),
    .p6(inst150_p6),
    .p7(inst150_p7),
    .p8(inst150_p8),
    .p9(inst150_p9),
    .reset(inst150_reset)
);
comp92 inst151 (
    .clk(inst151_clk),
    .p10(inst151_p10),
    .p11(inst151_p11),
    .p12(inst151_p12),
    .p13(inst151_p13),
    .p14(inst151_p14),
    .p15(inst151_p15),
    .p16(inst151_p16),
    .p17(inst151_p17),
    .p18(inst151_p18),
    .p19(inst151_p19),
    .p20(inst151_p20),
    .p21(inst151_p21),
    .p22(inst151_p22),
    .p23(inst151_p23),
    .p24(inst151_p24),
    .p25(inst151_p25),
    .p26(inst151_p26),
    .p27(inst151_p27),
    .p28(inst151_p28),
    .p29(inst151_p29),
    .p30(inst151_p30),
    .p31(inst151_p31),
    .p32(inst151_p32),
    .p33(inst151_p33),
    .p34(inst151_p34),
    .p35(inst151_p35),
    .p36(inst151_p36),
    .p37(inst151_p37),
    .p5(inst151_p5),
    .p6(inst151_p6),
    .p7(inst151_p7),
    .p8(inst151_p8),
    .p9(inst151_p9),
    .reset(inst151_reset)
);
comp93 inst152 (
    .clk(inst152_clk),
    .p10(inst152_p10),
    .p11(inst152_p11),
    .p12(inst152_p12),
    .p13(inst152_p13),
    .p14(inst152_p14),
    .p15(inst152_p15),
    .p16(inst152_p16),
    .p17(inst152_p17),
    .p18(inst152_p18),
    .p19(inst152_p19),
    .p20(inst152_p20),
    .p21(inst152_p21),
    .p22(inst152_p22),
    .p23(inst152_p23),
    .p24(inst152_p24),
    .p25(inst152_p25),
    .p26(inst152_p26),
    .p27(inst152_p27),
    .p28(inst152_p28),
    .p29(inst152_p29),
    .p30(inst152_p30),
    .p31(inst152_p31),
    .p32(inst152_p32),
    .p33(inst152_p33),
    .p34(inst152_p34),
    .p35(inst152_p35),
    .p36(inst152_p36),
    .p4(inst152_p4),
    .p5(inst152_p5),
    .p6(inst152_p6),
    .p7(inst152_p7),
    .p8(inst152_p8),
    .p9(inst152_p9),
    .reset(inst152_reset)
);
wire _guard0 = 1;
wire _guard1 = ev00__0state >= 6'd2;
wire _guard2 = ev00__0state <= 6'd2;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = ev00__0state >= 6'd41;
wire _guard5 = ev00__0state <= 6'd41;
wire _guard6 = _guard4 & _guard5;
wire _guard7 = ev00__0state >= 6'd31;
wire _guard8 = ev00__0state <= 6'd31;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = ev00__0state >= 6'd26;
wire _guard11 = ev00__0state <= 6'd26;
wire _guard12 = _guard10 & _guard11;
wire _guard13 = ev00__0state >= 6'd26;
wire _guard14 = ev00__0state <= 6'd26;
wire _guard15 = _guard13 & _guard14;
wire _guard16 = ev00__0state >= 6'd26;
wire _guard17 = ev00__0state <= 6'd26;
wire _guard18 = _guard16 & _guard17;
wire _guard19 = ev00__0state >= 6'd26;
wire _guard20 = ev00__0state <= 6'd26;
wire _guard21 = _guard19 & _guard20;
wire _guard22 = ev00__0state >= 6'd50;
wire _guard23 = ev00__0state <= 6'd50;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = ev00__0state >= 6'd50;
wire _guard26 = ev00__0state <= 6'd50;
wire _guard27 = _guard25 & _guard26;
wire _guard28 = ev00__0state >= 6'd50;
wire _guard29 = ev00__0state <= 6'd50;
wire _guard30 = _guard28 & _guard29;
wire _guard31 = ev00__0state >= 6'd50;
wire _guard32 = ev00__0state <= 6'd50;
wire _guard33 = _guard31 & _guard32;
wire _guard34 = ev00__0state >= 6'd51;
wire _guard35 = ev00__0state <= 6'd51;
wire _guard36 = _guard34 & _guard35;
wire _guard37 = ev00__0state >= 6'd51;
wire _guard38 = ev00__0state <= 6'd51;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = ev00__0state >= 6'd51;
wire _guard41 = ev00__0state <= 6'd51;
wire _guard42 = _guard40 & _guard41;
wire _guard43 = ev00__0state >= 6'd51;
wire _guard44 = ev00__0state <= 6'd51;
wire _guard45 = _guard43 & _guard44;
wire _guard46 = ev00__0state >= 6'd51;
wire _guard47 = ev00__0state <= 6'd51;
wire _guard48 = _guard46 & _guard47;
wire _guard49 = ev00__0state >= 6'd51;
wire _guard50 = ev00__0state <= 6'd51;
wire _guard51 = _guard49 & _guard50;
wire _guard52 = ev00__0state >= 6'd51;
wire _guard53 = ev00__0state <= 6'd51;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = ev00__0state >= 6'd51;
wire _guard56 = ev00__0state <= 6'd51;
wire _guard57 = _guard55 & _guard56;
wire _guard58 = ev00__0state >= 6'd51;
wire _guard59 = ev00__0state <= 6'd51;
wire _guard60 = _guard58 & _guard59;
wire _guard61 = ev00__0state >= 6'd51;
wire _guard62 = ev00__0state <= 6'd51;
wire _guard63 = _guard61 & _guard62;
wire _guard64 = ev00__0state >= 6'd51;
wire _guard65 = ev00__0state <= 6'd51;
wire _guard66 = _guard64 & _guard65;
wire _guard67 = ev00__0state >= 6'd51;
wire _guard68 = ev00__0state <= 6'd51;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = ev00__0state >= 6'd51;
wire _guard71 = ev00__0state <= 6'd51;
wire _guard72 = _guard70 & _guard71;
wire _guard73 = ev00__0state >= 6'd51;
wire _guard74 = ev00__0state <= 6'd51;
wire _guard75 = _guard73 & _guard74;
wire _guard76 = ev00__0state >= 6'd51;
wire _guard77 = ev00__0state <= 6'd51;
wire _guard78 = _guard76 & _guard77;
wire _guard79 = ev00__0state >= 6'd51;
wire _guard80 = ev00__0state <= 6'd51;
wire _guard81 = _guard79 & _guard80;
wire _guard82 = ev00__0state >= 6'd51;
wire _guard83 = ev00__0state <= 6'd51;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = ev00__0state >= 6'd51;
wire _guard86 = ev00__0state <= 6'd51;
wire _guard87 = _guard85 & _guard86;
wire _guard88 = ev00__0state >= 6'd51;
wire _guard89 = ev00__0state <= 6'd51;
wire _guard90 = _guard88 & _guard89;
wire _guard91 = ev00__0state >= 6'd51;
wire _guard92 = ev00__0state <= 6'd51;
wire _guard93 = _guard91 & _guard92;
wire _guard94 = ev00__0state >= 6'd51;
wire _guard95 = ev00__0state <= 6'd51;
wire _guard96 = _guard94 & _guard95;
wire _guard97 = ev00__0state >= 6'd51;
wire _guard98 = ev00__0state <= 6'd51;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = ev00__0state >= 6'd51;
wire _guard101 = ev00__0state <= 6'd51;
wire _guard102 = _guard100 & _guard101;
wire _guard103 = ev00__0state >= 6'd51;
wire _guard104 = ev00__0state <= 6'd51;
wire _guard105 = _guard103 & _guard104;
wire _guard106 = ev00__0state >= 6'd51;
wire _guard107 = ev00__0state <= 6'd51;
wire _guard108 = _guard106 & _guard107;
wire _guard109 = ev00__0state >= 6'd51;
wire _guard110 = ev00__0state <= 6'd51;
wire _guard111 = _guard109 & _guard110;
wire _guard112 = ev00__0state >= 6'd51;
wire _guard113 = ev00__0state <= 6'd51;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = ev00__0state >= 6'd51;
wire _guard116 = ev00__0state <= 6'd51;
wire _guard117 = _guard115 & _guard116;
wire _guard118 = ev00__0state >= 6'd51;
wire _guard119 = ev00__0state <= 6'd51;
wire _guard120 = _guard118 & _guard119;
wire _guard121 = ev00__0state >= 6'd51;
wire _guard122 = ev00__0state <= 6'd51;
wire _guard123 = _guard121 & _guard122;
wire _guard124 = ev00__0state >= 6'd51;
wire _guard125 = ev00__0state <= 6'd51;
wire _guard126 = _guard124 & _guard125;
wire _guard127 = ev00__0state >= 6'd51;
wire _guard128 = ev00__0state <= 6'd51;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = ev00__1_0;
wire _guard131 = ev00__1state >= 6'd1;
wire _guard132 = ev00__1state <= 6'd0;
wire _guard133 = _guard131 & _guard132;
wire _guard134 = _guard130 | _guard133;
wire _guard135 = ev00__1_0;
wire _guard136 = ev00__1state >= 6'd1;
wire _guard137 = ev00__1state <= 6'd0;
wire _guard138 = _guard136 & _guard137;
wire _guard139 = _guard135 | _guard138;
wire _guard140 = ev00__1_0;
wire _guard141 = ev00__1state >= 6'd1;
wire _guard142 = ev00__1state <= 6'd0;
wire _guard143 = _guard141 & _guard142;
wire _guard144 = _guard140 | _guard143;
wire _guard145 = ev00__1_0;
wire _guard146 = ev00__1state >= 6'd1;
wire _guard147 = ev00__1state <= 6'd0;
wire _guard148 = _guard146 & _guard147;
wire _guard149 = _guard145 | _guard148;
wire _guard150 = ev00__1_0;
wire _guard151 = ev00__1state >= 6'd1;
wire _guard152 = ev00__1state <= 6'd0;
wire _guard153 = _guard151 & _guard152;
wire _guard154 = _guard150 | _guard153;
wire _guard155 = ev00__1_0;
wire _guard156 = ev00__1state >= 6'd1;
wire _guard157 = ev00__1state <= 6'd0;
wire _guard158 = _guard156 & _guard157;
wire _guard159 = _guard155 | _guard158;
wire _guard160 = ev00__1_0;
wire _guard161 = ev00__1state >= 6'd1;
wire _guard162 = ev00__1state <= 6'd0;
wire _guard163 = _guard161 & _guard162;
wire _guard164 = _guard160 | _guard163;
wire _guard165 = ev00__1_0;
wire _guard166 = ev00__1state >= 6'd1;
wire _guard167 = ev00__1state <= 6'd0;
wire _guard168 = _guard166 & _guard167;
wire _guard169 = _guard165 | _guard168;
wire _guard170 = ev00__1_0;
wire _guard171 = ev00__1state >= 6'd1;
wire _guard172 = ev00__1state <= 6'd0;
wire _guard173 = _guard171 & _guard172;
wire _guard174 = _guard170 | _guard173;
wire _guard175 = ev00__1_0;
wire _guard176 = ev00__1state >= 6'd1;
wire _guard177 = ev00__1state <= 6'd0;
wire _guard178 = _guard176 & _guard177;
wire _guard179 = _guard175 | _guard178;
wire _guard180 = ev00__1_0;
wire _guard181 = ev00__1state >= 6'd1;
wire _guard182 = ev00__1state <= 6'd0;
wire _guard183 = _guard181 & _guard182;
wire _guard184 = _guard180 | _guard183;
wire _guard185 = ev00__1_0;
wire _guard186 = ev00__1state >= 6'd1;
wire _guard187 = ev00__1state <= 6'd0;
wire _guard188 = _guard186 & _guard187;
wire _guard189 = _guard185 | _guard188;
wire _guard190 = ev00__1_0;
wire _guard191 = ev00__1state >= 6'd1;
wire _guard192 = ev00__1state <= 6'd0;
wire _guard193 = _guard191 & _guard192;
wire _guard194 = _guard190 | _guard193;
wire _guard195 = ev00__1_0;
wire _guard196 = ev00__1state >= 6'd1;
wire _guard197 = ev00__1state <= 6'd0;
wire _guard198 = _guard196 & _guard197;
wire _guard199 = _guard195 | _guard198;
wire _guard200 = ev00__1_0;
wire _guard201 = ev00__1state >= 6'd1;
wire _guard202 = ev00__1state <= 6'd0;
wire _guard203 = _guard201 & _guard202;
wire _guard204 = _guard200 | _guard203;
wire _guard205 = ev00__1_0;
wire _guard206 = ev00__1state >= 6'd1;
wire _guard207 = ev00__1state <= 6'd0;
wire _guard208 = _guard206 & _guard207;
wire _guard209 = _guard205 | _guard208;
wire _guard210 = ev00__1_0;
wire _guard211 = ev00__1state >= 6'd1;
wire _guard212 = ev00__1state <= 6'd0;
wire _guard213 = _guard211 & _guard212;
wire _guard214 = _guard210 | _guard213;
wire _guard215 = ev00__1_0;
wire _guard216 = ev00__1state >= 6'd1;
wire _guard217 = ev00__1state <= 6'd0;
wire _guard218 = _guard216 & _guard217;
wire _guard219 = _guard215 | _guard218;
wire _guard220 = ev00__1_0;
wire _guard221 = ev00__1state >= 6'd1;
wire _guard222 = ev00__1state <= 6'd0;
wire _guard223 = _guard221 & _guard222;
wire _guard224 = _guard220 | _guard223;
wire _guard225 = ev00__1_0;
wire _guard226 = ev00__1state >= 6'd1;
wire _guard227 = ev00__1state <= 6'd0;
wire _guard228 = _guard226 & _guard227;
wire _guard229 = _guard225 | _guard228;
wire _guard230 = ev00__1_0;
wire _guard231 = ev00__1state >= 6'd1;
wire _guard232 = ev00__1state <= 6'd0;
wire _guard233 = _guard231 & _guard232;
wire _guard234 = _guard230 | _guard233;
wire _guard235 = ev00__1_0;
wire _guard236 = ev00__1state >= 6'd1;
wire _guard237 = ev00__1state <= 6'd0;
wire _guard238 = _guard236 & _guard237;
wire _guard239 = _guard235 | _guard238;
wire _guard240 = ev00__1_0;
wire _guard241 = ev00__1state >= 6'd1;
wire _guard242 = ev00__1state <= 6'd0;
wire _guard243 = _guard241 & _guard242;
wire _guard244 = _guard240 | _guard243;
wire _guard245 = ev00__1_0;
wire _guard246 = ev00__1state >= 6'd1;
wire _guard247 = ev00__1state <= 6'd0;
wire _guard248 = _guard246 & _guard247;
wire _guard249 = _guard245 | _guard248;
wire _guard250 = ev00__1_0;
wire _guard251 = ev00__1state >= 6'd1;
wire _guard252 = ev00__1state <= 6'd0;
wire _guard253 = _guard251 & _guard252;
wire _guard254 = _guard250 | _guard253;
wire _guard255 = ev00__1_0;
wire _guard256 = ev00__1state >= 6'd1;
wire _guard257 = ev00__1state <= 6'd0;
wire _guard258 = _guard256 & _guard257;
wire _guard259 = _guard255 | _guard258;
wire _guard260 = ev00__1_0;
wire _guard261 = ev00__1state >= 6'd1;
wire _guard262 = ev00__1state <= 6'd0;
wire _guard263 = _guard261 & _guard262;
wire _guard264 = _guard260 | _guard263;
wire _guard265 = ev00__1_0;
wire _guard266 = ev00__1state >= 6'd1;
wire _guard267 = ev00__1state <= 6'd0;
wire _guard268 = _guard266 & _guard267;
wire _guard269 = _guard265 | _guard268;
wire _guard270 = ev00__1_0;
wire _guard271 = ev00__1state >= 6'd1;
wire _guard272 = ev00__1state <= 6'd0;
wire _guard273 = _guard271 & _guard272;
wire _guard274 = _guard270 | _guard273;
wire _guard275 = ev00__1_0;
wire _guard276 = ev00__1state >= 6'd1;
wire _guard277 = ev00__1state <= 6'd0;
wire _guard278 = _guard276 & _guard277;
wire _guard279 = _guard275 | _guard278;
wire _guard280 = ev00__1_0;
wire _guard281 = ev00__1state >= 6'd1;
wire _guard282 = ev00__1state <= 6'd0;
wire _guard283 = _guard281 & _guard282;
wire _guard284 = _guard280 | _guard283;
wire _guard285 = ev00__1_0;
wire _guard286 = ev00__1state >= 6'd1;
wire _guard287 = ev00__1state <= 6'd0;
wire _guard288 = _guard286 & _guard287;
wire _guard289 = _guard285 | _guard288;
wire _guard290 = ev00__0state >= 6'd38;
wire _guard291 = ev00__0state <= 6'd38;
wire _guard292 = _guard290 & _guard291;
wire _guard293 = ev00__0state >= 6'd44;
wire _guard294 = ev00__0state <= 6'd44;
wire _guard295 = _guard293 & _guard294;
wire _guard296 = ev00__0state >= 6'd44;
wire _guard297 = ev00__0state <= 6'd44;
wire _guard298 = _guard296 & _guard297;
wire _guard299 = ev00__0state >= 6'd44;
wire _guard300 = ev00__0state <= 6'd44;
wire _guard301 = _guard299 & _guard300;
wire _guard302 = ev00__0state >= 6'd44;
wire _guard303 = ev00__0state <= 6'd44;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = ev00__0state >= 6'd13;
wire _guard306 = ev00__0state <= 6'd13;
wire _guard307 = _guard305 & _guard306;
wire _guard308 = ev00__0state >= 6'd13;
wire _guard309 = ev00__0state <= 6'd13;
wire _guard310 = _guard308 & _guard309;
wire _guard311 = ev00__0state >= 6'd13;
wire _guard312 = ev00__0state <= 6'd13;
wire _guard313 = _guard311 & _guard312;
wire _guard314 = ev00__0state >= 6'd13;
wire _guard315 = ev00__0state <= 6'd13;
wire _guard316 = _guard314 & _guard315;
wire _guard317 = ev00__0state >= 6'd19;
wire _guard318 = ev00__0state <= 6'd19;
wire _guard319 = _guard317 & _guard318;
wire _guard320 = ev00__0state >= 6'd19;
wire _guard321 = ev00__0state <= 6'd19;
wire _guard322 = _guard320 & _guard321;
wire _guard323 = ev00__0state >= 6'd19;
wire _guard324 = ev00__0state <= 6'd19;
wire _guard325 = _guard323 & _guard324;
wire _guard326 = ev00__0state >= 6'd19;
wire _guard327 = ev00__0state <= 6'd19;
wire _guard328 = _guard326 & _guard327;
wire _guard329 = ev00__0state >= 6'd33;
wire _guard330 = ev00__0state <= 6'd33;
wire _guard331 = _guard329 & _guard330;
wire _guard332 = ev00__0state >= 6'd33;
wire _guard333 = ev00__0state <= 6'd33;
wire _guard334 = _guard332 & _guard333;
wire _guard335 = ev00__0state >= 6'd33;
wire _guard336 = ev00__0state <= 6'd33;
wire _guard337 = _guard335 & _guard336;
wire _guard338 = ev00__0state >= 6'd33;
wire _guard339 = ev00__0state <= 6'd33;
wire _guard340 = _guard338 & _guard339;
wire _guard341 = ev00__0state >= 6'd38;
wire _guard342 = ev00__0state <= 6'd38;
wire _guard343 = _guard341 & _guard342;
wire _guard344 = ev00__0state >= 6'd39;
wire _guard345 = ev00__0state <= 6'd39;
wire _guard346 = _guard344 & _guard345;
wire _guard347 = ev00__0state >= 6'd39;
wire _guard348 = ev00__0state <= 6'd39;
wire _guard349 = _guard347 & _guard348;
wire _guard350 = ev00__0state >= 6'd39;
wire _guard351 = ev00__0state <= 6'd39;
wire _guard352 = _guard350 & _guard351;
wire _guard353 = ev00__0state >= 6'd39;
wire _guard354 = ev00__0state <= 6'd39;
wire _guard355 = _guard353 & _guard354;
wire _guard356 = ev00__0state >= 6'd43;
wire _guard357 = ev00__0state <= 6'd43;
wire _guard358 = _guard356 & _guard357;
wire _guard359 = ev00__0state >= 6'd13;
wire _guard360 = ev00__0state <= 6'd13;
wire _guard361 = _guard359 & _guard360;
wire _guard362 = ev00__0state >= 6'd13;
wire _guard363 = ev00__0state <= 6'd13;
wire _guard364 = _guard362 & _guard363;
wire _guard365 = ev00__0state >= 6'd13;
wire _guard366 = ev00__0state <= 6'd13;
wire _guard367 = _guard365 & _guard366;
wire _guard368 = ev00__0state >= 6'd13;
wire _guard369 = ev00__0state <= 6'd13;
wire _guard370 = _guard368 & _guard369;
wire _guard371 = ev00__0state >= 6'd23;
wire _guard372 = ev00__0state <= 6'd23;
wire _guard373 = _guard371 & _guard372;
wire _guard374 = ev00__0state >= 6'd23;
wire _guard375 = ev00__0state <= 6'd23;
wire _guard376 = _guard374 & _guard375;
wire _guard377 = ev00__0state >= 6'd23;
wire _guard378 = ev00__0state <= 6'd23;
wire _guard379 = _guard377 & _guard378;
wire _guard380 = ev00__0state >= 6'd23;
wire _guard381 = ev00__0state <= 6'd23;
wire _guard382 = _guard380 & _guard381;
wire _guard383 = ev00__0_0;
wire _guard384 = ev00__0state >= 6'd1;
wire _guard385 = ev00__0state <= 6'd51;
wire _guard386 = _guard384 & _guard385;
wire _guard387 = _guard383 | _guard386;
wire _guard388 = ev00__0_0;
wire _guard389 = ev00__0state >= 6'd1;
wire _guard390 = ev00__0state <= 6'd51;
wire _guard391 = _guard389 & _guard390;
wire _guard392 = _guard388 | _guard391;
wire _guard393 = ev00__0_0;
wire _guard394 = ev00__0state >= 6'd1;
wire _guard395 = ev00__0state <= 6'd51;
wire _guard396 = _guard394 & _guard395;
wire _guard397 = _guard393 | _guard396;
wire _guard398 = ev00__0_0;
wire _guard399 = ev00__0state >= 6'd1;
wire _guard400 = ev00__0state <= 6'd51;
wire _guard401 = _guard399 & _guard400;
wire _guard402 = _guard398 | _guard401;
wire _guard403 = ev00__0_0;
wire _guard404 = ev00__0state >= 6'd1;
wire _guard405 = ev00__0state <= 6'd51;
wire _guard406 = _guard404 & _guard405;
wire _guard407 = _guard403 | _guard406;
wire _guard408 = ev00__0_0;
wire _guard409 = ev00__0state >= 6'd1;
wire _guard410 = ev00__0state <= 6'd51;
wire _guard411 = _guard409 & _guard410;
wire _guard412 = _guard408 | _guard411;
wire _guard413 = ev00__0_0;
wire _guard414 = ev00__0state >= 6'd1;
wire _guard415 = ev00__0state <= 6'd51;
wire _guard416 = _guard414 & _guard415;
wire _guard417 = _guard413 | _guard416;
wire _guard418 = ev00__0_0;
wire _guard419 = ev00__0state >= 6'd1;
wire _guard420 = ev00__0state <= 6'd51;
wire _guard421 = _guard419 & _guard420;
wire _guard422 = _guard418 | _guard421;
wire _guard423 = ev00__0_0;
wire _guard424 = ev00__0state >= 6'd1;
wire _guard425 = ev00__0state <= 6'd51;
wire _guard426 = _guard424 & _guard425;
wire _guard427 = _guard423 | _guard426;
wire _guard428 = ev00__0_0;
wire _guard429 = ev00__0state >= 6'd1;
wire _guard430 = ev00__0state <= 6'd51;
wire _guard431 = _guard429 & _guard430;
wire _guard432 = _guard428 | _guard431;
wire _guard433 = ev00__0_0;
wire _guard434 = ev00__0state >= 6'd1;
wire _guard435 = ev00__0state <= 6'd51;
wire _guard436 = _guard434 & _guard435;
wire _guard437 = _guard433 | _guard436;
wire _guard438 = ev00__0_0;
wire _guard439 = ev00__0state >= 6'd1;
wire _guard440 = ev00__0state <= 6'd51;
wire _guard441 = _guard439 & _guard440;
wire _guard442 = _guard438 | _guard441;
wire _guard443 = ev00__0_0;
wire _guard444 = ev00__0state >= 6'd1;
wire _guard445 = ev00__0state <= 6'd51;
wire _guard446 = _guard444 & _guard445;
wire _guard447 = _guard443 | _guard446;
wire _guard448 = ev00__0_0;
wire _guard449 = ev00__0state >= 6'd1;
wire _guard450 = ev00__0state <= 6'd51;
wire _guard451 = _guard449 & _guard450;
wire _guard452 = _guard448 | _guard451;
wire _guard453 = ev00__0_0;
wire _guard454 = ev00__0state >= 6'd1;
wire _guard455 = ev00__0state <= 6'd51;
wire _guard456 = _guard454 & _guard455;
wire _guard457 = _guard453 | _guard456;
wire _guard458 = ev00__0_0;
wire _guard459 = ev00__0state >= 6'd1;
wire _guard460 = ev00__0state <= 6'd51;
wire _guard461 = _guard459 & _guard460;
wire _guard462 = _guard458 | _guard461;
wire _guard463 = ev00__0state >= 6'd38;
wire _guard464 = ev00__0state <= 6'd38;
wire _guard465 = _guard463 & _guard464;
wire _guard466 = ev00__0state >= 6'd25;
wire _guard467 = ev00__0state <= 6'd25;
wire _guard468 = _guard466 & _guard467;
wire _guard469 = ev00__0state >= 6'd26;
wire _guard470 = ev00__0state <= 6'd26;
wire _guard471 = _guard469 & _guard470;
wire _guard472 = ev00__0state >= 6'd26;
wire _guard473 = ev00__0state <= 6'd26;
wire _guard474 = _guard472 & _guard473;
wire _guard475 = ev00__0state >= 6'd26;
wire _guard476 = ev00__0state <= 6'd26;
wire _guard477 = _guard475 & _guard476;
wire _guard478 = ev00__0state >= 6'd26;
wire _guard479 = ev00__0state <= 6'd26;
wire _guard480 = _guard478 & _guard479;
wire _guard481 = ev00__0state >= 6'd38;
wire _guard482 = ev00__0state <= 6'd38;
wire _guard483 = _guard481 & _guard482;
wire _guard484 = ev00__0state >= 6'd46;
wire _guard485 = ev00__0state <= 6'd46;
wire _guard486 = _guard484 & _guard485;
wire _guard487 = ev00__0state >= 6'd46;
wire _guard488 = ev00__0state <= 6'd46;
wire _guard489 = _guard487 & _guard488;
wire _guard490 = ev00__0state >= 6'd46;
wire _guard491 = ev00__0state <= 6'd46;
wire _guard492 = _guard490 & _guard491;
wire _guard493 = ev00__0state >= 6'd46;
wire _guard494 = ev00__0state <= 6'd46;
wire _guard495 = _guard493 & _guard494;
wire _guard496 = ev00__0state >= 6'd22;
wire _guard497 = ev00__0state <= 6'd22;
wire _guard498 = _guard496 & _guard497;
wire _guard499 = ev00__0state >= 6'd22;
wire _guard500 = ev00__0state <= 6'd22;
wire _guard501 = _guard499 & _guard500;
wire _guard502 = ev00__0state >= 6'd22;
wire _guard503 = ev00__0state <= 6'd22;
wire _guard504 = _guard502 & _guard503;
wire _guard505 = ev00__0state >= 6'd22;
wire _guard506 = ev00__0state <= 6'd22;
wire _guard507 = _guard505 & _guard506;
wire _guard508 = ev00__0state >= 6'd38;
wire _guard509 = ev00__0state <= 6'd38;
wire _guard510 = _guard508 & _guard509;
wire _guard511 = ev00__0state >= 6'd13;
wire _guard512 = ev00__0state <= 6'd13;
wire _guard513 = _guard511 & _guard512;
wire _guard514 = ev00__0state >= 6'd13;
wire _guard515 = ev00__0state <= 6'd13;
wire _guard516 = _guard514 & _guard515;
wire _guard517 = ev00__0state >= 6'd13;
wire _guard518 = ev00__0state <= 6'd13;
wire _guard519 = _guard517 & _guard518;
wire _guard520 = ev00__0state >= 6'd13;
wire _guard521 = ev00__0state <= 6'd13;
wire _guard522 = _guard520 & _guard521;
wire _guard523 = ev00__0state >= 6'd17;
wire _guard524 = ev00__0state <= 6'd17;
wire _guard525 = _guard523 & _guard524;
wire _guard526 = ev00__0state >= 6'd17;
wire _guard527 = ev00__0state <= 6'd17;
wire _guard528 = _guard526 & _guard527;
wire _guard529 = ev00__0state >= 6'd17;
wire _guard530 = ev00__0state <= 6'd17;
wire _guard531 = _guard529 & _guard530;
wire _guard532 = ev00__0state >= 6'd17;
wire _guard533 = ev00__0state <= 6'd17;
wire _guard534 = _guard532 & _guard533;
wire _guard535 = ev00__0state >= 6'd27;
wire _guard536 = ev00__0state <= 6'd27;
wire _guard537 = _guard535 & _guard536;
wire _guard538 = ev00__0state >= 6'd3;
wire _guard539 = ev00__0state <= 6'd3;
wire _guard540 = _guard538 & _guard539;
wire _guard541 = ev00__0state >= 6'd13;
wire _guard542 = ev00__0state <= 6'd13;
wire _guard543 = _guard541 & _guard542;
wire _guard544 = ev00__0state >= 6'd13;
wire _guard545 = ev00__0state <= 6'd13;
wire _guard546 = _guard544 & _guard545;
wire _guard547 = ev00__0state >= 6'd13;
wire _guard548 = ev00__0state <= 6'd13;
wire _guard549 = _guard547 & _guard548;
wire _guard550 = ev00__0state >= 6'd13;
wire _guard551 = ev00__0state <= 6'd13;
wire _guard552 = _guard550 & _guard551;
wire _guard553 = ev00__0state >= 6'd25;
wire _guard554 = ev00__0state <= 6'd25;
wire _guard555 = _guard553 & _guard554;
wire _guard556 = ev00__0state >= 6'd26;
wire _guard557 = ev00__0state <= 6'd26;
wire _guard558 = _guard556 & _guard557;
wire _guard559 = ev00__0state >= 6'd26;
wire _guard560 = ev00__0state <= 6'd26;
wire _guard561 = _guard559 & _guard560;
wire _guard562 = ev00__0state >= 6'd26;
wire _guard563 = ev00__0state <= 6'd26;
wire _guard564 = _guard562 & _guard563;
wire _guard565 = ev00__0state >= 6'd26;
wire _guard566 = ev00__0state <= 6'd26;
wire _guard567 = _guard565 & _guard566;
wire _guard568 = ev00__0state >= 6'd33;
wire _guard569 = ev00__0state <= 6'd33;
wire _guard570 = _guard568 & _guard569;
wire _guard571 = ev00__0state >= 6'd12;
wire _guard572 = ev00__0state <= 6'd12;
wire _guard573 = _guard571 & _guard572;
wire _guard574 = ev00__0state >= 6'd12;
wire _guard575 = ev00__0state <= 6'd12;
wire _guard576 = _guard574 & _guard575;
wire _guard577 = ev00__0state >= 6'd12;
wire _guard578 = ev00__0state <= 6'd12;
wire _guard579 = _guard577 & _guard578;
wire _guard580 = ev00__0state >= 6'd12;
wire _guard581 = ev00__0state <= 6'd12;
wire _guard582 = _guard580 & _guard581;
wire _guard583 = ev00__0state >= 6'd12;
wire _guard584 = ev00__0state <= 6'd12;
wire _guard585 = _guard583 & _guard584;
wire _guard586 = ev00__0state >= 6'd12;
wire _guard587 = ev00__0state <= 6'd12;
wire _guard588 = _guard586 & _guard587;
wire _guard589 = ev00__0state >= 6'd12;
wire _guard590 = ev00__0state <= 6'd12;
wire _guard591 = _guard589 & _guard590;
wire _guard592 = ev00__0state >= 6'd12;
wire _guard593 = ev00__0state <= 6'd12;
wire _guard594 = _guard592 & _guard593;
wire _guard595 = ev00__0state >= 6'd12;
wire _guard596 = ev00__0state <= 6'd12;
wire _guard597 = _guard595 & _guard596;
wire _guard598 = ev00__0state >= 6'd12;
wire _guard599 = ev00__0state <= 6'd12;
wire _guard600 = _guard598 & _guard599;
wire _guard601 = ev00__0state >= 6'd12;
wire _guard602 = ev00__0state <= 6'd12;
wire _guard603 = _guard601 & _guard602;
wire _guard604 = ev00__0state >= 6'd12;
wire _guard605 = ev00__0state <= 6'd12;
wire _guard606 = _guard604 & _guard605;
wire _guard607 = ev00__0state >= 6'd12;
wire _guard608 = ev00__0state <= 6'd12;
wire _guard609 = _guard607 & _guard608;
wire _guard610 = ev00__0state >= 6'd12;
wire _guard611 = ev00__0state <= 6'd12;
wire _guard612 = _guard610 & _guard611;
wire _guard613 = ev00__0state >= 6'd12;
wire _guard614 = ev00__0state <= 6'd12;
wire _guard615 = _guard613 & _guard614;
wire _guard616 = ev00__0state >= 6'd12;
wire _guard617 = ev00__0state <= 6'd12;
wire _guard618 = _guard616 & _guard617;
wire _guard619 = ev00__0state >= 6'd12;
wire _guard620 = ev00__0state <= 6'd12;
wire _guard621 = _guard619 & _guard620;
wire _guard622 = ev00__0state >= 6'd12;
wire _guard623 = ev00__0state <= 6'd12;
wire _guard624 = _guard622 & _guard623;
wire _guard625 = ev00__0state >= 6'd12;
wire _guard626 = ev00__0state <= 6'd12;
wire _guard627 = _guard625 & _guard626;
wire _guard628 = ev00__0state >= 6'd12;
wire _guard629 = ev00__0state <= 6'd12;
wire _guard630 = _guard628 & _guard629;
wire _guard631 = ev00__0state >= 6'd12;
wire _guard632 = ev00__0state <= 6'd12;
wire _guard633 = _guard631 & _guard632;
wire _guard634 = ev00__0state >= 6'd12;
wire _guard635 = ev00__0state <= 6'd12;
wire _guard636 = _guard634 & _guard635;
wire _guard637 = ev00__0state >= 6'd12;
wire _guard638 = ev00__0state <= 6'd12;
wire _guard639 = _guard637 & _guard638;
wire _guard640 = ev00__0state >= 6'd12;
wire _guard641 = ev00__0state <= 6'd12;
wire _guard642 = _guard640 & _guard641;
wire _guard643 = ev00__0state >= 6'd12;
wire _guard644 = ev00__0state <= 6'd12;
wire _guard645 = _guard643 & _guard644;
wire _guard646 = ev00__0state >= 6'd12;
wire _guard647 = ev00__0state <= 6'd12;
wire _guard648 = _guard646 & _guard647;
wire _guard649 = ev00__0state >= 6'd12;
wire _guard650 = ev00__0state <= 6'd12;
wire _guard651 = _guard649 & _guard650;
wire _guard652 = ev00__0state >= 6'd12;
wire _guard653 = ev00__0state <= 6'd12;
wire _guard654 = _guard652 & _guard653;
wire _guard655 = ev00__0state >= 6'd12;
wire _guard656 = ev00__0state <= 6'd12;
wire _guard657 = _guard655 & _guard656;
wire _guard658 = ev00__0state >= 6'd12;
wire _guard659 = ev00__0state <= 6'd12;
wire _guard660 = _guard658 & _guard659;
wire _guard661 = ev00__0state >= 6'd12;
wire _guard662 = ev00__0state <= 6'd12;
wire _guard663 = _guard661 & _guard662;
wire _guard664 = ev00__0state >= 6'd12;
wire _guard665 = ev00__0state <= 6'd12;
wire _guard666 = _guard664 & _guard665;
wire _guard667 = ev00__0_0;
wire _guard668 = ev00__0state >= 6'd1;
wire _guard669 = ev00__0state <= 6'd51;
wire _guard670 = _guard668 & _guard669;
wire _guard671 = _guard667 | _guard670;
wire _guard672 = ev00__0_0;
wire _guard673 = ev00__0state >= 6'd1;
wire _guard674 = ev00__0state <= 6'd51;
wire _guard675 = _guard673 & _guard674;
wire _guard676 = _guard672 | _guard675;
wire _guard677 = ev00__0_0;
wire _guard678 = ev00__0state >= 6'd1;
wire _guard679 = ev00__0state <= 6'd51;
wire _guard680 = _guard678 & _guard679;
wire _guard681 = _guard677 | _guard680;
wire _guard682 = ev00__0_0;
wire _guard683 = ev00__0state >= 6'd1;
wire _guard684 = ev00__0state <= 6'd51;
wire _guard685 = _guard683 & _guard684;
wire _guard686 = _guard682 | _guard685;
wire _guard687 = ev00__0_0;
wire _guard688 = ev00__0state >= 6'd1;
wire _guard689 = ev00__0state <= 6'd51;
wire _guard690 = _guard688 & _guard689;
wire _guard691 = _guard687 | _guard690;
wire _guard692 = ev00__0_0;
wire _guard693 = ev00__0state >= 6'd1;
wire _guard694 = ev00__0state <= 6'd51;
wire _guard695 = _guard693 & _guard694;
wire _guard696 = _guard692 | _guard695;
wire _guard697 = ev00__0_0;
wire _guard698 = ev00__0state >= 6'd1;
wire _guard699 = ev00__0state <= 6'd51;
wire _guard700 = _guard698 & _guard699;
wire _guard701 = _guard697 | _guard700;
wire _guard702 = ev00__0_0;
wire _guard703 = ev00__0state >= 6'd1;
wire _guard704 = ev00__0state <= 6'd51;
wire _guard705 = _guard703 & _guard704;
wire _guard706 = _guard702 | _guard705;
wire _guard707 = ev00__0_0;
wire _guard708 = ev00__0state >= 6'd1;
wire _guard709 = ev00__0state <= 6'd51;
wire _guard710 = _guard708 & _guard709;
wire _guard711 = _guard707 | _guard710;
wire _guard712 = ev00__0_0;
wire _guard713 = ev00__0state >= 6'd1;
wire _guard714 = ev00__0state <= 6'd51;
wire _guard715 = _guard713 & _guard714;
wire _guard716 = _guard712 | _guard715;
wire _guard717 = ev00__0_0;
wire _guard718 = ev00__0state >= 6'd1;
wire _guard719 = ev00__0state <= 6'd51;
wire _guard720 = _guard718 & _guard719;
wire _guard721 = _guard717 | _guard720;
wire _guard722 = ev00__0_0;
wire _guard723 = ev00__0state >= 6'd1;
wire _guard724 = ev00__0state <= 6'd51;
wire _guard725 = _guard723 & _guard724;
wire _guard726 = _guard722 | _guard725;
wire _guard727 = ev00__0_0;
wire _guard728 = ev00__0state >= 6'd1;
wire _guard729 = ev00__0state <= 6'd51;
wire _guard730 = _guard728 & _guard729;
wire _guard731 = _guard727 | _guard730;
wire _guard732 = ev00__0_0;
wire _guard733 = ev00__0state >= 6'd1;
wire _guard734 = ev00__0state <= 6'd51;
wire _guard735 = _guard733 & _guard734;
wire _guard736 = _guard732 | _guard735;
wire _guard737 = ev00__0_0;
wire _guard738 = ev00__0state >= 6'd1;
wire _guard739 = ev00__0state <= 6'd51;
wire _guard740 = _guard738 & _guard739;
wire _guard741 = _guard737 | _guard740;
wire _guard742 = ev00__0_0;
wire _guard743 = ev00__0state >= 6'd1;
wire _guard744 = ev00__0state <= 6'd51;
wire _guard745 = _guard743 & _guard744;
wire _guard746 = _guard742 | _guard745;
wire _guard747 = ev00__0state >= 6'd4;
wire _guard748 = ev00__0state <= 6'd4;
wire _guard749 = _guard747 & _guard748;
wire _guard750 = ev00__0state >= 6'd4;
wire _guard751 = ev00__0state <= 6'd4;
wire _guard752 = _guard750 & _guard751;
wire _guard753 = ev00__0state >= 6'd4;
wire _guard754 = ev00__0state <= 6'd4;
wire _guard755 = _guard753 & _guard754;
wire _guard756 = ev00__0state >= 6'd4;
wire _guard757 = ev00__0state <= 6'd4;
wire _guard758 = _guard756 & _guard757;
wire _guard759 = ev00__0state >= 6'd14;
wire _guard760 = ev00__0state <= 6'd14;
wire _guard761 = _guard759 & _guard760;
wire _guard762 = ev00__0state >= 6'd13;
wire _guard763 = ev00__0state <= 6'd13;
wire _guard764 = _guard762 & _guard763;
wire _guard765 = ev00__0state >= 6'd13;
wire _guard766 = ev00__0state <= 6'd13;
wire _guard767 = _guard765 & _guard766;
wire _guard768 = ev00__0state >= 6'd13;
wire _guard769 = ev00__0state <= 6'd13;
wire _guard770 = _guard768 & _guard769;
wire _guard771 = ev00__0state >= 6'd13;
wire _guard772 = ev00__0state <= 6'd13;
wire _guard773 = _guard771 & _guard772;
wire _guard774 = ev00__0state >= 6'd25;
wire _guard775 = ev00__0state <= 6'd25;
wire _guard776 = _guard774 & _guard775;
wire _guard777 = ev00__0state >= 6'd9;
wire _guard778 = ev00__0state <= 6'd9;
wire _guard779 = _guard777 & _guard778;
wire _guard780 = ev00__0state >= 6'd9;
wire _guard781 = ev00__0state <= 6'd9;
wire _guard782 = _guard780 & _guard781;
wire _guard783 = ev00__0state >= 6'd9;
wire _guard784 = ev00__0state <= 6'd9;
wire _guard785 = _guard783 & _guard784;
wire _guard786 = ev00__0state >= 6'd9;
wire _guard787 = ev00__0state <= 6'd9;
wire _guard788 = _guard786 & _guard787;
wire _guard789 = ev00__0state >= 6'd38;
wire _guard790 = ev00__0state <= 6'd38;
wire _guard791 = _guard789 & _guard790;
wire _guard792 = ev00__0state >= 6'd39;
wire _guard793 = ev00__0state <= 6'd39;
wire _guard794 = _guard792 & _guard793;
wire _guard795 = ev00__0state >= 6'd39;
wire _guard796 = ev00__0state <= 6'd39;
wire _guard797 = _guard795 & _guard796;
wire _guard798 = ev00__0state >= 6'd39;
wire _guard799 = ev00__0state <= 6'd39;
wire _guard800 = _guard798 & _guard799;
wire _guard801 = ev00__0state >= 6'd39;
wire _guard802 = ev00__0state <= 6'd39;
wire _guard803 = _guard801 & _guard802;
wire _guard804 = ev00__0state >= 6'd32;
wire _guard805 = ev00__0state <= 6'd32;
wire _guard806 = _guard804 & _guard805;
wire _guard807 = ev00__1_0;
wire _guard808 = ev00__1state >= 6'd1;
wire _guard809 = ev00__1state <= 6'd0;
wire _guard810 = _guard808 & _guard809;
wire _guard811 = _guard807 | _guard810;
wire _guard812 = ev00__0_0;
wire _guard813 = ev00__0state >= 6'd1;
wire _guard814 = ev00__0state <= 6'd0;
wire _guard815 = _guard813 & _guard814;
wire _guard816 = _guard812 | _guard815;
wire _guard817 = ev00__0_0;
wire _guard818 = ev00__0state >= 6'd1;
wire _guard819 = ev00__0state <= 6'd0;
wire _guard820 = _guard818 & _guard819;
wire _guard821 = _guard817 | _guard820;
wire _guard822 = ev00__0_0;
wire _guard823 = ev00__0state >= 6'd1;
wire _guard824 = ev00__0state <= 6'd0;
wire _guard825 = _guard823 & _guard824;
wire _guard826 = _guard822 | _guard825;
wire _guard827 = ev00__0_0;
wire _guard828 = ev00__0state >= 6'd1;
wire _guard829 = ev00__0state <= 6'd0;
wire _guard830 = _guard828 & _guard829;
wire _guard831 = _guard827 | _guard830;
wire _guard832 = ev00__0_0;
wire _guard833 = ev00__0state >= 6'd1;
wire _guard834 = ev00__0state <= 6'd0;
wire _guard835 = _guard833 & _guard834;
wire _guard836 = _guard832 | _guard835;
wire _guard837 = ev00__0_0;
wire _guard838 = ev00__0state >= 6'd1;
wire _guard839 = ev00__0state <= 6'd0;
wire _guard840 = _guard838 & _guard839;
wire _guard841 = _guard837 | _guard840;
wire _guard842 = ev00__0_0;
wire _guard843 = ev00__0state >= 6'd1;
wire _guard844 = ev00__0state <= 6'd0;
wire _guard845 = _guard843 & _guard844;
wire _guard846 = _guard842 | _guard845;
wire _guard847 = ev00__0_0;
wire _guard848 = ev00__0state >= 6'd1;
wire _guard849 = ev00__0state <= 6'd0;
wire _guard850 = _guard848 & _guard849;
wire _guard851 = _guard847 | _guard850;
wire _guard852 = ev00__0_0;
wire _guard853 = ev00__0state >= 6'd1;
wire _guard854 = ev00__0state <= 6'd0;
wire _guard855 = _guard853 & _guard854;
wire _guard856 = _guard852 | _guard855;
wire _guard857 = ev00__0_0;
wire _guard858 = ev00__0state >= 6'd1;
wire _guard859 = ev00__0state <= 6'd0;
wire _guard860 = _guard858 & _guard859;
wire _guard861 = _guard857 | _guard860;
wire _guard862 = ev00__0_0;
wire _guard863 = ev00__0state >= 6'd1;
wire _guard864 = ev00__0state <= 6'd0;
wire _guard865 = _guard863 & _guard864;
wire _guard866 = _guard862 | _guard865;
wire _guard867 = ev00__0_0;
wire _guard868 = ev00__0state >= 6'd1;
wire _guard869 = ev00__0state <= 6'd0;
wire _guard870 = _guard868 & _guard869;
wire _guard871 = _guard867 | _guard870;
wire _guard872 = ev00__0_0;
wire _guard873 = ev00__0state >= 6'd1;
wire _guard874 = ev00__0state <= 6'd0;
wire _guard875 = _guard873 & _guard874;
wire _guard876 = _guard872 | _guard875;
wire _guard877 = ev00__0_0;
wire _guard878 = ev00__0state >= 6'd1;
wire _guard879 = ev00__0state <= 6'd0;
wire _guard880 = _guard878 & _guard879;
wire _guard881 = _guard877 | _guard880;
wire _guard882 = ev00__0_0;
wire _guard883 = ev00__0state >= 6'd1;
wire _guard884 = ev00__0state <= 6'd0;
wire _guard885 = _guard883 & _guard884;
wire _guard886 = _guard882 | _guard885;
wire _guard887 = ev00__0_0;
wire _guard888 = ev00__0state >= 6'd1;
wire _guard889 = ev00__0state <= 6'd0;
wire _guard890 = _guard888 & _guard889;
wire _guard891 = _guard887 | _guard890;
wire _guard892 = ev00__0_0;
wire _guard893 = ev00__0state >= 6'd1;
wire _guard894 = ev00__0state <= 6'd0;
wire _guard895 = _guard893 & _guard894;
wire _guard896 = _guard892 | _guard895;
wire _guard897 = ev00__0_0;
wire _guard898 = ev00__0state >= 6'd1;
wire _guard899 = ev00__0state <= 6'd0;
wire _guard900 = _guard898 & _guard899;
wire _guard901 = _guard897 | _guard900;
wire _guard902 = ev00__0_0;
wire _guard903 = ev00__0state >= 6'd1;
wire _guard904 = ev00__0state <= 6'd0;
wire _guard905 = _guard903 & _guard904;
wire _guard906 = _guard902 | _guard905;
wire _guard907 = ev00__0_0;
wire _guard908 = ev00__0state >= 6'd1;
wire _guard909 = ev00__0state <= 6'd0;
wire _guard910 = _guard908 & _guard909;
wire _guard911 = _guard907 | _guard910;
wire _guard912 = ev00__0_0;
wire _guard913 = ev00__0state >= 6'd1;
wire _guard914 = ev00__0state <= 6'd0;
wire _guard915 = _guard913 & _guard914;
wire _guard916 = _guard912 | _guard915;
wire _guard917 = ev00__0_0;
wire _guard918 = ev00__0state >= 6'd1;
wire _guard919 = ev00__0state <= 6'd0;
wire _guard920 = _guard918 & _guard919;
wire _guard921 = _guard917 | _guard920;
wire _guard922 = ev00__0_0;
wire _guard923 = ev00__0state >= 6'd1;
wire _guard924 = ev00__0state <= 6'd0;
wire _guard925 = _guard923 & _guard924;
wire _guard926 = _guard922 | _guard925;
wire _guard927 = ev00__0_0;
wire _guard928 = ev00__0state >= 6'd1;
wire _guard929 = ev00__0state <= 6'd0;
wire _guard930 = _guard928 & _guard929;
wire _guard931 = _guard927 | _guard930;
wire _guard932 = ev00__0_0;
wire _guard933 = ev00__0state >= 6'd1;
wire _guard934 = ev00__0state <= 6'd0;
wire _guard935 = _guard933 & _guard934;
wire _guard936 = _guard932 | _guard935;
wire _guard937 = ev00__0_0;
wire _guard938 = ev00__0state >= 6'd1;
wire _guard939 = ev00__0state <= 6'd0;
wire _guard940 = _guard938 & _guard939;
wire _guard941 = _guard937 | _guard940;
wire _guard942 = ev00__0_0;
wire _guard943 = ev00__0state >= 6'd1;
wire _guard944 = ev00__0state <= 6'd0;
wire _guard945 = _guard943 & _guard944;
wire _guard946 = _guard942 | _guard945;
wire _guard947 = ev00__0_0;
wire _guard948 = ev00__0state >= 6'd1;
wire _guard949 = ev00__0state <= 6'd0;
wire _guard950 = _guard948 & _guard949;
wire _guard951 = _guard947 | _guard950;
wire _guard952 = ev00__0_0;
wire _guard953 = ev00__0state >= 6'd1;
wire _guard954 = ev00__0state <= 6'd0;
wire _guard955 = _guard953 & _guard954;
wire _guard956 = _guard952 | _guard955;
wire _guard957 = ev00__0_0;
wire _guard958 = ev00__0state >= 6'd1;
wire _guard959 = ev00__0state <= 6'd0;
wire _guard960 = _guard958 & _guard959;
wire _guard961 = _guard957 | _guard960;
wire _guard962 = ev00__0_0;
wire _guard963 = ev00__0state >= 6'd1;
wire _guard964 = ev00__0state <= 6'd0;
wire _guard965 = _guard963 & _guard964;
wire _guard966 = _guard962 | _guard965;
wire _guard967 = ev00__0_0;
wire _guard968 = ev00__0state >= 6'd1;
wire _guard969 = ev00__0state <= 6'd0;
wire _guard970 = _guard968 & _guard969;
wire _guard971 = _guard967 | _guard970;
wire _guard972 = ev00__0state >= 6'd51;
wire _guard973 = ev00__0state <= 6'd51;
wire _guard974 = _guard972 & _guard973;
wire _guard975 = ev00__0state >= 6'd5;
wire _guard976 = ev00__0state <= 6'd5;
wire _guard977 = _guard975 & _guard976;
wire _guard978 = ev00__0state >= 6'd5;
wire _guard979 = ev00__0state <= 6'd5;
wire _guard980 = _guard978 & _guard979;
wire _guard981 = ev00__0state >= 6'd5;
wire _guard982 = ev00__0state <= 6'd5;
wire _guard983 = _guard981 & _guard982;
wire _guard984 = ev00__0state >= 6'd5;
wire _guard985 = ev00__0state <= 6'd5;
wire _guard986 = _guard984 & _guard985;
wire _guard987 = ev00__0_0;
wire _guard988 = ev00__0state >= 6'd1;
wire _guard989 = ev00__0state <= 6'd0;
wire _guard990 = _guard988 & _guard989;
wire _guard991 = _guard987 | _guard990;
wire _guard992 = ev00__0state >= 6'd6;
wire _guard993 = ev00__0state <= 6'd6;
wire _guard994 = _guard992 & _guard993;
wire _guard995 = _guard991 | _guard994;
wire _guard996 = ev00__0state >= 6'd13;
wire _guard997 = ev00__0state <= 6'd13;
wire _guard998 = _guard996 & _guard997;
wire _guard999 = _guard995 | _guard998;
wire _guard1000 = ev00__0state >= 6'd19;
wire _guard1001 = ev00__0state <= 6'd19;
wire _guard1002 = _guard1000 & _guard1001;
wire _guard1003 = _guard999 | _guard1002;
wire _guard1004 = ev00__0state >= 6'd26;
wire _guard1005 = ev00__0state <= 6'd26;
wire _guard1006 = _guard1004 & _guard1005;
wire _guard1007 = _guard1003 | _guard1006;
wire _guard1008 = ev00__0state >= 6'd32;
wire _guard1009 = ev00__0state <= 6'd32;
wire _guard1010 = _guard1008 & _guard1009;
wire _guard1011 = _guard1007 | _guard1010;
wire _guard1012 = ev00__0state >= 6'd39;
wire _guard1013 = ev00__0state <= 6'd39;
wire _guard1014 = _guard1012 & _guard1013;
wire _guard1015 = _guard1011 | _guard1014;
wire _guard1016 = ev00__0state >= 6'd45;
wire _guard1017 = ev00__0state <= 6'd45;
wire _guard1018 = _guard1016 & _guard1017;
wire _guard1019 = _guard1015 | _guard1018;
wire _guard1020 = ev00__0state >= 6'd13;
wire _guard1021 = ev00__0state <= 6'd13;
wire _guard1022 = _guard1020 & _guard1021;
wire _guard1023 = ev00__0state >= 6'd19;
wire _guard1024 = ev00__0state <= 6'd19;
wire _guard1025 = _guard1023 & _guard1024;
wire _guard1026 = ev00__0state >= 6'd26;
wire _guard1027 = ev00__0state <= 6'd26;
wire _guard1028 = _guard1026 & _guard1027;
wire _guard1029 = ev00__0state >= 6'd45;
wire _guard1030 = ev00__0state <= 6'd45;
wire _guard1031 = _guard1029 & _guard1030;
wire _guard1032 = ev00__0state >= 6'd39;
wire _guard1033 = ev00__0state <= 6'd39;
wire _guard1034 = _guard1032 & _guard1033;
wire _guard1035 = ev00__0state >= 6'd32;
wire _guard1036 = ev00__0state <= 6'd32;
wire _guard1037 = _guard1035 & _guard1036;
wire _guard1038 = ev00__0_0;
wire _guard1039 = ev00__0state >= 6'd1;
wire _guard1040 = ev00__0state <= 6'd0;
wire _guard1041 = _guard1039 & _guard1040;
wire _guard1042 = _guard1038 | _guard1041;
wire _guard1043 = ev00__0state >= 6'd6;
wire _guard1044 = ev00__0state <= 6'd6;
wire _guard1045 = _guard1043 & _guard1044;
wire _guard1046 = ev00__0_0;
wire _guard1047 = ev00__0state >= 6'd1;
wire _guard1048 = ev00__0state <= 6'd0;
wire _guard1049 = _guard1047 & _guard1048;
wire _guard1050 = _guard1046 | _guard1049;
wire _guard1051 = ev00__0state >= 6'd9;
wire _guard1052 = ev00__0state <= 6'd9;
wire _guard1053 = _guard1051 & _guard1052;
wire _guard1054 = _guard1050 | _guard1053;
wire _guard1055 = ev00__0state >= 6'd13;
wire _guard1056 = ev00__0state <= 6'd13;
wire _guard1057 = _guard1055 & _guard1056;
wire _guard1058 = _guard1054 | _guard1057;
wire _guard1059 = ev00__0state >= 6'd22;
wire _guard1060 = ev00__0state <= 6'd22;
wire _guard1061 = _guard1059 & _guard1060;
wire _guard1062 = _guard1058 | _guard1061;
wire _guard1063 = ev00__0state >= 6'd26;
wire _guard1064 = ev00__0state <= 6'd26;
wire _guard1065 = _guard1063 & _guard1064;
wire _guard1066 = _guard1062 | _guard1065;
wire _guard1067 = ev00__0state >= 6'd35;
wire _guard1068 = ev00__0state <= 6'd35;
wire _guard1069 = _guard1067 & _guard1068;
wire _guard1070 = _guard1066 | _guard1069;
wire _guard1071 = ev00__0state >= 6'd39;
wire _guard1072 = ev00__0state <= 6'd39;
wire _guard1073 = _guard1071 & _guard1072;
wire _guard1074 = _guard1070 | _guard1073;
wire _guard1075 = ev00__0state >= 6'd48;
wire _guard1076 = ev00__0state <= 6'd48;
wire _guard1077 = _guard1075 & _guard1076;
wire _guard1078 = _guard1074 | _guard1077;
wire _guard1079 = ev00__0state >= 6'd22;
wire _guard1080 = ev00__0state <= 6'd22;
wire _guard1081 = _guard1079 & _guard1080;
wire _guard1082 = ev00__0state >= 6'd26;
wire _guard1083 = ev00__0state <= 6'd26;
wire _guard1084 = _guard1082 & _guard1083;
wire _guard1085 = ev00__0state >= 6'd9;
wire _guard1086 = ev00__0state <= 6'd9;
wire _guard1087 = _guard1085 & _guard1086;
wire _guard1088 = ev00__0state >= 6'd39;
wire _guard1089 = ev00__0state <= 6'd39;
wire _guard1090 = _guard1088 & _guard1089;
wire _guard1091 = ev00__0state >= 6'd13;
wire _guard1092 = ev00__0state <= 6'd13;
wire _guard1093 = _guard1091 & _guard1092;
wire _guard1094 = ev00__0state >= 6'd48;
wire _guard1095 = ev00__0state <= 6'd48;
wire _guard1096 = _guard1094 & _guard1095;
wire _guard1097 = ev00__0_0;
wire _guard1098 = ev00__0state >= 6'd1;
wire _guard1099 = ev00__0state <= 6'd0;
wire _guard1100 = _guard1098 & _guard1099;
wire _guard1101 = _guard1097 | _guard1100;
wire _guard1102 = ev00__0state >= 6'd35;
wire _guard1103 = ev00__0state <= 6'd35;
wire _guard1104 = _guard1102 & _guard1103;
wire _guard1105 = ev00__0state >= 6'd5;
wire _guard1106 = ev00__0state <= 6'd5;
wire _guard1107 = _guard1105 & _guard1106;
wire _guard1108 = ev00__0_0;
wire _guard1109 = ev00__0state >= 6'd1;
wire _guard1110 = ev00__0state <= 6'd0;
wire _guard1111 = _guard1109 & _guard1110;
wire _guard1112 = _guard1108 | _guard1111;
wire _guard1113 = ev00__0state >= 6'd10;
wire _guard1114 = ev00__0state <= 6'd10;
wire _guard1115 = _guard1113 & _guard1114;
wire _guard1116 = _guard1112 | _guard1115;
wire _guard1117 = ev00__0state >= 6'd13;
wire _guard1118 = ev00__0state <= 6'd13;
wire _guard1119 = _guard1117 & _guard1118;
wire _guard1120 = _guard1116 | _guard1119;
wire _guard1121 = ev00__0state >= 6'd23;
wire _guard1122 = ev00__0state <= 6'd23;
wire _guard1123 = _guard1121 & _guard1122;
wire _guard1124 = _guard1120 | _guard1123;
wire _guard1125 = ev00__0state >= 6'd26;
wire _guard1126 = ev00__0state <= 6'd26;
wire _guard1127 = _guard1125 & _guard1126;
wire _guard1128 = _guard1124 | _guard1127;
wire _guard1129 = ev00__0state >= 6'd36;
wire _guard1130 = ev00__0state <= 6'd36;
wire _guard1131 = _guard1129 & _guard1130;
wire _guard1132 = _guard1128 | _guard1131;
wire _guard1133 = ev00__0state >= 6'd39;
wire _guard1134 = ev00__0state <= 6'd39;
wire _guard1135 = _guard1133 & _guard1134;
wire _guard1136 = _guard1132 | _guard1135;
wire _guard1137 = ev00__0state >= 6'd49;
wire _guard1138 = ev00__0state <= 6'd49;
wire _guard1139 = _guard1137 & _guard1138;
wire _guard1140 = _guard1136 | _guard1139;
wire _guard1141 = ev00__0state >= 6'd13;
wire _guard1142 = ev00__0state <= 6'd13;
wire _guard1143 = _guard1141 & _guard1142;
wire _guard1144 = ev00__0state >= 6'd23;
wire _guard1145 = ev00__0state <= 6'd23;
wire _guard1146 = _guard1144 & _guard1145;
wire _guard1147 = ev00__0state >= 6'd39;
wire _guard1148 = ev00__0state <= 6'd39;
wire _guard1149 = _guard1147 & _guard1148;
wire _guard1150 = ev00__0state >= 6'd10;
wire _guard1151 = ev00__0state <= 6'd10;
wire _guard1152 = _guard1150 & _guard1151;
wire _guard1153 = ev00__0state >= 6'd49;
wire _guard1154 = ev00__0state <= 6'd49;
wire _guard1155 = _guard1153 & _guard1154;
wire _guard1156 = ev00__0state >= 6'd26;
wire _guard1157 = ev00__0state <= 6'd26;
wire _guard1158 = _guard1156 & _guard1157;
wire _guard1159 = ev00__0_0;
wire _guard1160 = ev00__0state >= 6'd1;
wire _guard1161 = ev00__0state <= 6'd0;
wire _guard1162 = _guard1160 & _guard1161;
wire _guard1163 = _guard1159 | _guard1162;
wire _guard1164 = ev00__0state >= 6'd36;
wire _guard1165 = ev00__0state <= 6'd36;
wire _guard1166 = _guard1164 & _guard1165;
wire _guard1167 = ev00__0state >= 6'd45;
wire _guard1168 = ev00__0state <= 6'd45;
wire _guard1169 = _guard1167 & _guard1168;
wire _guard1170 = ev00__0state >= 6'd39;
wire _guard1171 = ev00__0state <= 6'd39;
wire _guard1172 = _guard1170 & _guard1171;
wire _guard1173 = ev00__0state >= 6'd39;
wire _guard1174 = ev00__0state <= 6'd39;
wire _guard1175 = _guard1173 & _guard1174;
wire _guard1176 = ev00__0state >= 6'd39;
wire _guard1177 = ev00__0state <= 6'd39;
wire _guard1178 = _guard1176 & _guard1177;
wire _guard1179 = ev00__0state >= 6'd39;
wire _guard1180 = ev00__0state <= 6'd39;
wire _guard1181 = _guard1179 & _guard1180;
wire _guard1182 = ev00__0state >= 6'd25;
wire _guard1183 = ev00__0state <= 6'd25;
wire _guard1184 = _guard1182 & _guard1183;
wire _guard1185 = ev00__0_0;
wire _guard1186 = ev00__0state >= 6'd1;
wire _guard1187 = ev00__0state <= 6'd0;
wire _guard1188 = _guard1186 & _guard1187;
wire _guard1189 = _guard1185 | _guard1188;
wire _guard1190 = ev00__0_0;
wire _guard1191 = ev00__0state >= 6'd1;
wire _guard1192 = ev00__0state <= 6'd0;
wire _guard1193 = _guard1191 & _guard1192;
wire _guard1194 = _guard1190 | _guard1193;
wire _guard1195 = ev00__0_0;
wire _guard1196 = ev00__0state >= 6'd1;
wire _guard1197 = ev00__0state <= 6'd0;
wire _guard1198 = _guard1196 & _guard1197;
wire _guard1199 = _guard1195 | _guard1198;
wire _guard1200 = ev00__0_0;
wire _guard1201 = ev00__0state >= 6'd1;
wire _guard1202 = ev00__0state <= 6'd0;
wire _guard1203 = _guard1201 & _guard1202;
wire _guard1204 = _guard1200 | _guard1203;
wire _guard1205 = ev00__0state >= 6'd40;
wire _guard1206 = ev00__0state <= 6'd40;
wire _guard1207 = _guard1205 & _guard1206;
wire _guard1208 = ev00__0state >= 6'd51;
wire _guard1209 = ev00__0state <= 6'd51;
wire _guard1210 = _guard1208 & _guard1209;
wire _guard1211 = ev00__0state >= 6'd25;
wire _guard1212 = ev00__0state <= 6'd25;
wire _guard1213 = _guard1211 & _guard1212;
wire _guard1214 = ev00__0state >= 6'd28;
wire _guard1215 = ev00__0state <= 6'd28;
wire _guard1216 = _guard1214 & _guard1215;
wire _guard1217 = ev00__0state >= 6'd51;
wire _guard1218 = ev00__0state <= 6'd51;
wire _guard1219 = _guard1217 & _guard1218;
wire _guard1220 = ev00__0state >= 6'd17;
wire _guard1221 = ev00__0state <= 6'd17;
wire _guard1222 = _guard1220 & _guard1221;
wire _guard1223 = ev00__0state >= 6'd26;
wire _guard1224 = ev00__0state <= 6'd26;
wire _guard1225 = _guard1223 & _guard1224;
wire _guard1226 = ev00__0state >= 6'd26;
wire _guard1227 = ev00__0state <= 6'd26;
wire _guard1228 = _guard1226 & _guard1227;
wire _guard1229 = ev00__0state >= 6'd26;
wire _guard1230 = ev00__0state <= 6'd26;
wire _guard1231 = _guard1229 & _guard1230;
wire _guard1232 = ev00__0state >= 6'd26;
wire _guard1233 = ev00__0state <= 6'd26;
wire _guard1234 = _guard1232 & _guard1233;
wire _guard1235 = ev00__0state >= 6'd19;
wire _guard1236 = ev00__0state <= 6'd19;
wire _guard1237 = _guard1235 & _guard1236;
wire _guard1238 = ev00__0state >= 6'd11;
wire _guard1239 = ev00__0state <= 6'd11;
wire _guard1240 = _guard1238 & _guard1239;
wire _guard1241 = ev00__0state >= 6'd11;
wire _guard1242 = ev00__0state <= 6'd11;
wire _guard1243 = _guard1241 & _guard1242;
wire _guard1244 = ev00__0state >= 6'd11;
wire _guard1245 = ev00__0state <= 6'd11;
wire _guard1246 = _guard1244 & _guard1245;
wire _guard1247 = ev00__0state >= 6'd11;
wire _guard1248 = ev00__0state <= 6'd11;
wire _guard1249 = _guard1247 & _guard1248;
wire _guard1250 = ev00__0state >= 6'd12;
wire _guard1251 = ev00__0state <= 6'd12;
wire _guard1252 = _guard1250 & _guard1251;
wire _guard1253 = ev00__0state >= 6'd13;
wire _guard1254 = ev00__0state <= 6'd13;
wire _guard1255 = _guard1253 & _guard1254;
wire _guard1256 = ev00__0state >= 6'd13;
wire _guard1257 = ev00__0state <= 6'd13;
wire _guard1258 = _guard1256 & _guard1257;
wire _guard1259 = ev00__0state >= 6'd13;
wire _guard1260 = ev00__0state <= 6'd13;
wire _guard1261 = _guard1259 & _guard1260;
wire _guard1262 = ev00__0state >= 6'd13;
wire _guard1263 = ev00__0state <= 6'd13;
wire _guard1264 = _guard1262 & _guard1263;
wire _guard1265 = ev00__0state >= 6'd37;
wire _guard1266 = ev00__0state <= 6'd37;
wire _guard1267 = _guard1265 & _guard1266;
wire _guard1268 = ev00__0state >= 6'd37;
wire _guard1269 = ev00__0state <= 6'd37;
wire _guard1270 = _guard1268 & _guard1269;
wire _guard1271 = ev00__0state >= 6'd37;
wire _guard1272 = ev00__0state <= 6'd37;
wire _guard1273 = _guard1271 & _guard1272;
wire _guard1274 = ev00__0state >= 6'd37;
wire _guard1275 = ev00__0state <= 6'd37;
wire _guard1276 = _guard1274 & _guard1275;
wire _guard1277 = ev00__0state >= 6'd25;
wire _guard1278 = ev00__0state <= 6'd25;
wire _guard1279 = _guard1277 & _guard1278;
wire _guard1280 = ev00__0state >= 6'd25;
wire _guard1281 = ev00__0state <= 6'd25;
wire _guard1282 = _guard1280 & _guard1281;
wire _guard1283 = ev00__0state >= 6'd25;
wire _guard1284 = ev00__0state <= 6'd25;
wire _guard1285 = _guard1283 & _guard1284;
wire _guard1286 = ev00__0state >= 6'd25;
wire _guard1287 = ev00__0state <= 6'd25;
wire _guard1288 = _guard1286 & _guard1287;
wire _guard1289 = ev00__0state >= 6'd25;
wire _guard1290 = ev00__0state <= 6'd25;
wire _guard1291 = _guard1289 & _guard1290;
wire _guard1292 = ev00__0state >= 6'd25;
wire _guard1293 = ev00__0state <= 6'd25;
wire _guard1294 = _guard1292 & _guard1293;
wire _guard1295 = ev00__0state >= 6'd25;
wire _guard1296 = ev00__0state <= 6'd25;
wire _guard1297 = _guard1295 & _guard1296;
wire _guard1298 = ev00__0state >= 6'd25;
wire _guard1299 = ev00__0state <= 6'd25;
wire _guard1300 = _guard1298 & _guard1299;
wire _guard1301 = ev00__0state >= 6'd25;
wire _guard1302 = ev00__0state <= 6'd25;
wire _guard1303 = _guard1301 & _guard1302;
wire _guard1304 = ev00__0state >= 6'd25;
wire _guard1305 = ev00__0state <= 6'd25;
wire _guard1306 = _guard1304 & _guard1305;
wire _guard1307 = ev00__0state >= 6'd25;
wire _guard1308 = ev00__0state <= 6'd25;
wire _guard1309 = _guard1307 & _guard1308;
wire _guard1310 = ev00__0state >= 6'd25;
wire _guard1311 = ev00__0state <= 6'd25;
wire _guard1312 = _guard1310 & _guard1311;
wire _guard1313 = ev00__0state >= 6'd25;
wire _guard1314 = ev00__0state <= 6'd25;
wire _guard1315 = _guard1313 & _guard1314;
wire _guard1316 = ev00__0state >= 6'd25;
wire _guard1317 = ev00__0state <= 6'd25;
wire _guard1318 = _guard1316 & _guard1317;
wire _guard1319 = ev00__0state >= 6'd25;
wire _guard1320 = ev00__0state <= 6'd25;
wire _guard1321 = _guard1319 & _guard1320;
wire _guard1322 = ev00__0state >= 6'd25;
wire _guard1323 = ev00__0state <= 6'd25;
wire _guard1324 = _guard1322 & _guard1323;
wire _guard1325 = ev00__0state >= 6'd25;
wire _guard1326 = ev00__0state <= 6'd25;
wire _guard1327 = _guard1325 & _guard1326;
wire _guard1328 = ev00__0state >= 6'd25;
wire _guard1329 = ev00__0state <= 6'd25;
wire _guard1330 = _guard1328 & _guard1329;
wire _guard1331 = ev00__0state >= 6'd25;
wire _guard1332 = ev00__0state <= 6'd25;
wire _guard1333 = _guard1331 & _guard1332;
wire _guard1334 = ev00__0state >= 6'd25;
wire _guard1335 = ev00__0state <= 6'd25;
wire _guard1336 = _guard1334 & _guard1335;
wire _guard1337 = ev00__0state >= 6'd25;
wire _guard1338 = ev00__0state <= 6'd25;
wire _guard1339 = _guard1337 & _guard1338;
wire _guard1340 = ev00__0state >= 6'd25;
wire _guard1341 = ev00__0state <= 6'd25;
wire _guard1342 = _guard1340 & _guard1341;
wire _guard1343 = ev00__0state >= 6'd25;
wire _guard1344 = ev00__0state <= 6'd25;
wire _guard1345 = _guard1343 & _guard1344;
wire _guard1346 = ev00__0state >= 6'd25;
wire _guard1347 = ev00__0state <= 6'd25;
wire _guard1348 = _guard1346 & _guard1347;
wire _guard1349 = ev00__0state >= 6'd25;
wire _guard1350 = ev00__0state <= 6'd25;
wire _guard1351 = _guard1349 & _guard1350;
wire _guard1352 = ev00__0state >= 6'd25;
wire _guard1353 = ev00__0state <= 6'd25;
wire _guard1354 = _guard1352 & _guard1353;
wire _guard1355 = ev00__0state >= 6'd25;
wire _guard1356 = ev00__0state <= 6'd25;
wire _guard1357 = _guard1355 & _guard1356;
wire _guard1358 = ev00__0state >= 6'd25;
wire _guard1359 = ev00__0state <= 6'd25;
wire _guard1360 = _guard1358 & _guard1359;
wire _guard1361 = ev00__0state >= 6'd25;
wire _guard1362 = ev00__0state <= 6'd25;
wire _guard1363 = _guard1361 & _guard1362;
wire _guard1364 = ev00__0state >= 6'd25;
wire _guard1365 = ev00__0state <= 6'd25;
wire _guard1366 = _guard1364 & _guard1365;
wire _guard1367 = ev00__0state >= 6'd25;
wire _guard1368 = ev00__0state <= 6'd25;
wire _guard1369 = _guard1367 & _guard1368;
wire _guard1370 = ev00__0state >= 6'd25;
wire _guard1371 = ev00__0state <= 6'd25;
wire _guard1372 = _guard1370 & _guard1371;
wire _guard1373 = ev00__0state >= 6'd26;
wire _guard1374 = ev00__0state <= 6'd26;
wire _guard1375 = _guard1373 & _guard1374;
wire _guard1376 = ev00__0_0;
wire _guard1377 = ev00__0state >= 6'd1;
wire _guard1378 = ev00__0state <= 6'd0;
wire _guard1379 = _guard1377 & _guard1378;
wire _guard1380 = _guard1376 | _guard1379;
wire _guard1381 = ev00__0state >= 6'd4;
wire _guard1382 = ev00__0state <= 6'd4;
wire _guard1383 = _guard1381 & _guard1382;
wire _guard1384 = _guard1380 | _guard1383;
wire _guard1385 = ev00__0state >= 6'd13;
wire _guard1386 = ev00__0state <= 6'd13;
wire _guard1387 = _guard1385 & _guard1386;
wire _guard1388 = _guard1384 | _guard1387;
wire _guard1389 = ev00__0state >= 6'd17;
wire _guard1390 = ev00__0state <= 6'd17;
wire _guard1391 = _guard1389 & _guard1390;
wire _guard1392 = _guard1388 | _guard1391;
wire _guard1393 = ev00__0state >= 6'd26;
wire _guard1394 = ev00__0state <= 6'd26;
wire _guard1395 = _guard1393 & _guard1394;
wire _guard1396 = _guard1392 | _guard1395;
wire _guard1397 = ev00__0state >= 6'd30;
wire _guard1398 = ev00__0state <= 6'd30;
wire _guard1399 = _guard1397 & _guard1398;
wire _guard1400 = _guard1396 | _guard1399;
wire _guard1401 = ev00__0state >= 6'd39;
wire _guard1402 = ev00__0state <= 6'd39;
wire _guard1403 = _guard1401 & _guard1402;
wire _guard1404 = _guard1400 | _guard1403;
wire _guard1405 = ev00__0state >= 6'd43;
wire _guard1406 = ev00__0state <= 6'd43;
wire _guard1407 = _guard1405 & _guard1406;
wire _guard1408 = _guard1404 | _guard1407;
wire _guard1409 = ev00__0state >= 6'd13;
wire _guard1410 = ev00__0state <= 6'd13;
wire _guard1411 = _guard1409 & _guard1410;
wire _guard1412 = ev00__0state >= 6'd17;
wire _guard1413 = ev00__0state <= 6'd17;
wire _guard1414 = _guard1412 & _guard1413;
wire _guard1415 = ev00__0state >= 6'd4;
wire _guard1416 = ev00__0state <= 6'd4;
wire _guard1417 = _guard1415 & _guard1416;
wire _guard1418 = ev00__0state >= 6'd43;
wire _guard1419 = ev00__0state <= 6'd43;
wire _guard1420 = _guard1418 & _guard1419;
wire _guard1421 = ev00__0state >= 6'd39;
wire _guard1422 = ev00__0state <= 6'd39;
wire _guard1423 = _guard1421 & _guard1422;
wire _guard1424 = ev00__0state >= 6'd26;
wire _guard1425 = ev00__0state <= 6'd26;
wire _guard1426 = _guard1424 & _guard1425;
wire _guard1427 = ev00__0state >= 6'd30;
wire _guard1428 = ev00__0state <= 6'd30;
wire _guard1429 = _guard1427 & _guard1428;
wire _guard1430 = ev00__0_0;
wire _guard1431 = ev00__0state >= 6'd1;
wire _guard1432 = ev00__0state <= 6'd0;
wire _guard1433 = _guard1431 & _guard1432;
wire _guard1434 = _guard1430 | _guard1433;
wire _guard1435 = ev00__0state >= 6'd25;
wire _guard1436 = ev00__0state <= 6'd25;
wire _guard1437 = _guard1435 & _guard1436;
wire _guard1438 = ev00__0state >= 6'd15;
wire _guard1439 = ev00__0state <= 6'd15;
wire _guard1440 = _guard1438 & _guard1439;
wire _guard1441 = ev00__0_0;
wire _guard1442 = ev00__0state >= 6'd1;
wire _guard1443 = ev00__0state <= 6'd0;
wire _guard1444 = _guard1442 & _guard1443;
wire _guard1445 = _guard1441 | _guard1444;
wire _guard1446 = ev00__0_0;
wire _guard1447 = ev00__0state >= 6'd1;
wire _guard1448 = ev00__0state <= 6'd0;
wire _guard1449 = _guard1447 & _guard1448;
wire _guard1450 = _guard1446 | _guard1449;
wire _guard1451 = ev00__0_0;
wire _guard1452 = ev00__0state >= 6'd1;
wire _guard1453 = ev00__0state <= 6'd0;
wire _guard1454 = _guard1452 & _guard1453;
wire _guard1455 = _guard1451 | _guard1454;
wire _guard1456 = ev00__0_0;
wire _guard1457 = ev00__0state >= 6'd1;
wire _guard1458 = ev00__0state <= 6'd0;
wire _guard1459 = _guard1457 & _guard1458;
wire _guard1460 = _guard1456 | _guard1459;
wire _guard1461 = ev00__0state >= 6'd26;
wire _guard1462 = ev00__0state <= 6'd26;
wire _guard1463 = _guard1461 & _guard1462;
wire _guard1464 = ev00__0state >= 6'd26;
wire _guard1465 = ev00__0state <= 6'd26;
wire _guard1466 = _guard1464 & _guard1465;
wire _guard1467 = ev00__0state >= 6'd26;
wire _guard1468 = ev00__0state <= 6'd26;
wire _guard1469 = _guard1467 & _guard1468;
wire _guard1470 = ev00__0state >= 6'd26;
wire _guard1471 = ev00__0state <= 6'd26;
wire _guard1472 = _guard1470 & _guard1471;
wire _guard1473 = ev00__0state >= 6'd51;
wire _guard1474 = ev00__0state <= 6'd51;
wire _guard1475 = _guard1473 & _guard1474;
wire _guard1476 = ev00__0state >= 6'd39;
wire _guard1477 = ev00__0state <= 6'd39;
wire _guard1478 = _guard1476 & _guard1477;
wire _guard1479 = ev00__0state >= 6'd43;
wire _guard1480 = ev00__0state <= 6'd43;
wire _guard1481 = _guard1479 & _guard1480;
wire _guard1482 = ev00__0state >= 6'd43;
wire _guard1483 = ev00__0state <= 6'd43;
wire _guard1484 = _guard1482 & _guard1483;
wire _guard1485 = ev00__0state >= 6'd43;
wire _guard1486 = ev00__0state <= 6'd43;
wire _guard1487 = _guard1485 & _guard1486;
wire _guard1488 = ev00__0state >= 6'd43;
wire _guard1489 = ev00__0state <= 6'd43;
wire _guard1490 = _guard1488 & _guard1489;
wire _guard1491 = ev00__0state >= 6'd45;
wire _guard1492 = ev00__0state <= 6'd45;
wire _guard1493 = _guard1491 & _guard1492;
wire _guard1494 = ev00__0state >= 6'd45;
wire _guard1495 = ev00__0state <= 6'd45;
wire _guard1496 = _guard1494 & _guard1495;
wire _guard1497 = ev00__0state >= 6'd45;
wire _guard1498 = ev00__0state <= 6'd45;
wire _guard1499 = _guard1497 & _guard1498;
wire _guard1500 = ev00__0state >= 6'd45;
wire _guard1501 = ev00__0state <= 6'd45;
wire _guard1502 = _guard1500 & _guard1501;
wire _guard1503 = ev00__0state >= 6'd4;
wire _guard1504 = ev00__0state <= 6'd4;
wire _guard1505 = _guard1503 & _guard1504;
wire _guard1506 = ev00__0state >= 6'd13;
wire _guard1507 = ev00__0state <= 6'd13;
wire _guard1508 = _guard1506 & _guard1507;
wire _guard1509 = ev00__0state >= 6'd13;
wire _guard1510 = ev00__0state <= 6'd13;
wire _guard1511 = _guard1509 & _guard1510;
wire _guard1512 = ev00__0state >= 6'd13;
wire _guard1513 = ev00__0state <= 6'd13;
wire _guard1514 = _guard1512 & _guard1513;
wire _guard1515 = ev00__0state >= 6'd13;
wire _guard1516 = ev00__0state <= 6'd13;
wire _guard1517 = _guard1515 & _guard1516;
wire _guard1518 = ev00__0_0;
wire _guard1519 = ev00__0state >= 6'd1;
wire _guard1520 = ev00__0state <= 6'd0;
wire _guard1521 = _guard1519 & _guard1520;
wire _guard1522 = _guard1518 | _guard1521;
wire _guard1523 = ev00__0state >= 6'd11;
wire _guard1524 = ev00__0state <= 6'd11;
wire _guard1525 = _guard1523 & _guard1524;
wire _guard1526 = _guard1522 | _guard1525;
wire _guard1527 = ev00__0state >= 6'd13;
wire _guard1528 = ev00__0state <= 6'd13;
wire _guard1529 = _guard1527 & _guard1528;
wire _guard1530 = _guard1526 | _guard1529;
wire _guard1531 = ev00__0state >= 6'd24;
wire _guard1532 = ev00__0state <= 6'd24;
wire _guard1533 = _guard1531 & _guard1532;
wire _guard1534 = _guard1530 | _guard1533;
wire _guard1535 = ev00__0state >= 6'd26;
wire _guard1536 = ev00__0state <= 6'd26;
wire _guard1537 = _guard1535 & _guard1536;
wire _guard1538 = _guard1534 | _guard1537;
wire _guard1539 = ev00__0state >= 6'd37;
wire _guard1540 = ev00__0state <= 6'd37;
wire _guard1541 = _guard1539 & _guard1540;
wire _guard1542 = _guard1538 | _guard1541;
wire _guard1543 = ev00__0state >= 6'd39;
wire _guard1544 = ev00__0state <= 6'd39;
wire _guard1545 = _guard1543 & _guard1544;
wire _guard1546 = _guard1542 | _guard1545;
wire _guard1547 = ev00__0state >= 6'd50;
wire _guard1548 = ev00__0state <= 6'd50;
wire _guard1549 = _guard1547 & _guard1548;
wire _guard1550 = _guard1546 | _guard1549;
wire _guard1551 = ev00__0state >= 6'd26;
wire _guard1552 = ev00__0state <= 6'd26;
wire _guard1553 = _guard1551 & _guard1552;
wire _guard1554 = ev00__0state >= 6'd50;
wire _guard1555 = ev00__0state <= 6'd50;
wire _guard1556 = _guard1554 & _guard1555;
wire _guard1557 = ev00__0state >= 6'd11;
wire _guard1558 = ev00__0state <= 6'd11;
wire _guard1559 = _guard1557 & _guard1558;
wire _guard1560 = ev00__0state >= 6'd13;
wire _guard1561 = ev00__0state <= 6'd13;
wire _guard1562 = _guard1560 & _guard1561;
wire _guard1563 = ev00__0state >= 6'd37;
wire _guard1564 = ev00__0state <= 6'd37;
wire _guard1565 = _guard1563 & _guard1564;
wire _guard1566 = ev00__0_0;
wire _guard1567 = ev00__0state >= 6'd1;
wire _guard1568 = ev00__0state <= 6'd0;
wire _guard1569 = _guard1567 & _guard1568;
wire _guard1570 = _guard1566 | _guard1569;
wire _guard1571 = ev00__0state >= 6'd24;
wire _guard1572 = ev00__0state <= 6'd24;
wire _guard1573 = _guard1571 & _guard1572;
wire _guard1574 = ev00__0state >= 6'd39;
wire _guard1575 = ev00__0state <= 6'd39;
wire _guard1576 = _guard1574 & _guard1575;
wire _guard1577 = ev00__0state >= 6'd46;
wire _guard1578 = ev00__0state <= 6'd46;
wire _guard1579 = _guard1577 & _guard1578;
wire _guard1580 = ev00__0state >= 6'd5;
wire _guard1581 = ev00__0state <= 6'd5;
wire _guard1582 = _guard1580 & _guard1581;
wire _guard1583 = ev00__0state >= 6'd1;
wire _guard1584 = ev00__0state <= 6'd1;
wire _guard1585 = _guard1583 & _guard1584;
wire _guard1586 = ev00__0_0;
wire _guard1587 = ev00__0state >= 6'd1;
wire _guard1588 = ev00__0state <= 6'd0;
wire _guard1589 = _guard1587 & _guard1588;
wire _guard1590 = _guard1586 | _guard1589;
wire _guard1591 = ev00__0state >= 6'd6;
wire _guard1592 = ev00__0state <= 6'd6;
wire _guard1593 = _guard1591 & _guard1592;
wire _guard1594 = ev00__0state >= 6'd3;
wire _guard1595 = ev00__0state <= 6'd3;
wire _guard1596 = _guard1594 & _guard1595;
wire _guard1597 = ev00__0state >= 6'd7;
wire _guard1598 = ev00__0state <= 6'd7;
wire _guard1599 = _guard1597 & _guard1598;
wire _guard1600 = ev00__0state >= 6'd4;
wire _guard1601 = ev00__0state <= 6'd4;
wire _guard1602 = _guard1600 & _guard1601;
wire _guard1603 = ev00__0state >= 6'd2;
wire _guard1604 = ev00__0state <= 6'd2;
wire _guard1605 = _guard1603 & _guard1604;
wire _guard1606 = ev00__0state >= 6'd44;
wire _guard1607 = ev00__0state <= 6'd44;
wire _guard1608 = _guard1606 & _guard1607;
wire _guard1609 = ev00__0state >= 6'd40;
wire _guard1610 = ev00__0state <= 6'd40;
wire _guard1611 = _guard1609 & _guard1610;
wire _guard1612 = ev00__0state >= 6'd39;
wire _guard1613 = ev00__0state <= 6'd39;
wire _guard1614 = _guard1612 & _guard1613;
wire _guard1615 = ev00__0state >= 6'd45;
wire _guard1616 = ev00__0state <= 6'd45;
wire _guard1617 = _guard1615 & _guard1616;
wire _guard1618 = ev00__0state >= 6'd42;
wire _guard1619 = ev00__0state <= 6'd42;
wire _guard1620 = _guard1618 & _guard1619;
wire _guard1621 = ev00__0state >= 6'd46;
wire _guard1622 = ev00__0state <= 6'd46;
wire _guard1623 = _guard1621 & _guard1622;
wire _guard1624 = ev00__0state >= 6'd43;
wire _guard1625 = ev00__0state <= 6'd43;
wire _guard1626 = _guard1624 & _guard1625;
wire _guard1627 = ev00__0state >= 6'd41;
wire _guard1628 = ev00__0state <= 6'd41;
wire _guard1629 = _guard1627 & _guard1628;
wire _guard1630 = ev00__0state >= 6'd31;
wire _guard1631 = ev00__0state <= 6'd31;
wire _guard1632 = _guard1630 & _guard1631;
wire _guard1633 = ev00__0state >= 6'd27;
wire _guard1634 = ev00__0state <= 6'd27;
wire _guard1635 = _guard1633 & _guard1634;
wire _guard1636 = ev00__0state >= 6'd26;
wire _guard1637 = ev00__0state <= 6'd26;
wire _guard1638 = _guard1636 & _guard1637;
wire _guard1639 = ev00__0state >= 6'd32;
wire _guard1640 = ev00__0state <= 6'd32;
wire _guard1641 = _guard1639 & _guard1640;
wire _guard1642 = ev00__0state >= 6'd29;
wire _guard1643 = ev00__0state <= 6'd29;
wire _guard1644 = _guard1642 & _guard1643;
wire _guard1645 = ev00__0state >= 6'd33;
wire _guard1646 = ev00__0state <= 6'd33;
wire _guard1647 = _guard1645 & _guard1646;
wire _guard1648 = ev00__0state >= 6'd30;
wire _guard1649 = ev00__0state <= 6'd30;
wire _guard1650 = _guard1648 & _guard1649;
wire _guard1651 = ev00__0state >= 6'd28;
wire _guard1652 = ev00__0state <= 6'd28;
wire _guard1653 = _guard1651 & _guard1652;
wire _guard1654 = ev00__0state >= 6'd18;
wire _guard1655 = ev00__0state <= 6'd18;
wire _guard1656 = _guard1654 & _guard1655;
wire _guard1657 = ev00__0state >= 6'd14;
wire _guard1658 = ev00__0state <= 6'd14;
wire _guard1659 = _guard1657 & _guard1658;
wire _guard1660 = ev00__0state >= 6'd13;
wire _guard1661 = ev00__0state <= 6'd13;
wire _guard1662 = _guard1660 & _guard1661;
wire _guard1663 = ev00__0state >= 6'd19;
wire _guard1664 = ev00__0state <= 6'd19;
wire _guard1665 = _guard1663 & _guard1664;
wire _guard1666 = ev00__0state >= 6'd16;
wire _guard1667 = ev00__0state <= 6'd16;
wire _guard1668 = _guard1666 & _guard1667;
wire _guard1669 = ev00__0state >= 6'd20;
wire _guard1670 = ev00__0state <= 6'd20;
wire _guard1671 = _guard1669 & _guard1670;
wire _guard1672 = ev00__0state >= 6'd17;
wire _guard1673 = ev00__0state <= 6'd17;
wire _guard1674 = _guard1672 & _guard1673;
wire _guard1675 = ev00__0state >= 6'd15;
wire _guard1676 = ev00__0state <= 6'd15;
wire _guard1677 = _guard1675 & _guard1676;
wire _guard1678 = ev00__0_0;
wire _guard1679 = ev00__0state >= 6'd1;
wire _guard1680 = ev00__0state <= 6'd0;
wire _guard1681 = _guard1679 & _guard1680;
wire _guard1682 = _guard1678 | _guard1681;
wire _guard1683 = ev00__0state >= 6'd13;
wire _guard1684 = ev00__0state <= 6'd13;
wire _guard1685 = _guard1683 & _guard1684;
wire _guard1686 = _guard1682 | _guard1685;
wire _guard1687 = ev00__0state >= 6'd26;
wire _guard1688 = ev00__0state <= 6'd26;
wire _guard1689 = _guard1687 & _guard1688;
wire _guard1690 = _guard1686 | _guard1689;
wire _guard1691 = ev00__0state >= 6'd39;
wire _guard1692 = ev00__0state <= 6'd39;
wire _guard1693 = _guard1691 & _guard1692;
wire _guard1694 = _guard1690 | _guard1693;
wire _guard1695 = ev00__0state >= 6'd1;
wire _guard1696 = ev00__0state <= 6'd1;
wire _guard1697 = _guard1695 & _guard1696;
wire _guard1698 = _guard1694 | _guard1697;
wire _guard1699 = ev00__0state >= 6'd14;
wire _guard1700 = ev00__0state <= 6'd14;
wire _guard1701 = _guard1699 & _guard1700;
wire _guard1702 = _guard1698 | _guard1701;
wire _guard1703 = ev00__0state >= 6'd27;
wire _guard1704 = ev00__0state <= 6'd27;
wire _guard1705 = _guard1703 & _guard1704;
wire _guard1706 = _guard1702 | _guard1705;
wire _guard1707 = ev00__0state >= 6'd40;
wire _guard1708 = ev00__0state <= 6'd40;
wire _guard1709 = _guard1707 & _guard1708;
wire _guard1710 = _guard1706 | _guard1709;
wire _guard1711 = ev00__0state >= 6'd2;
wire _guard1712 = ev00__0state <= 6'd2;
wire _guard1713 = _guard1711 & _guard1712;
wire _guard1714 = _guard1710 | _guard1713;
wire _guard1715 = ev00__0state >= 6'd15;
wire _guard1716 = ev00__0state <= 6'd15;
wire _guard1717 = _guard1715 & _guard1716;
wire _guard1718 = _guard1714 | _guard1717;
wire _guard1719 = ev00__0state >= 6'd28;
wire _guard1720 = ev00__0state <= 6'd28;
wire _guard1721 = _guard1719 & _guard1720;
wire _guard1722 = _guard1718 | _guard1721;
wire _guard1723 = ev00__0state >= 6'd41;
wire _guard1724 = ev00__0state <= 6'd41;
wire _guard1725 = _guard1723 & _guard1724;
wire _guard1726 = _guard1722 | _guard1725;
wire _guard1727 = ev00__0state >= 6'd3;
wire _guard1728 = ev00__0state <= 6'd3;
wire _guard1729 = _guard1727 & _guard1728;
wire _guard1730 = _guard1726 | _guard1729;
wire _guard1731 = ev00__0state >= 6'd16;
wire _guard1732 = ev00__0state <= 6'd16;
wire _guard1733 = _guard1731 & _guard1732;
wire _guard1734 = _guard1730 | _guard1733;
wire _guard1735 = ev00__0state >= 6'd29;
wire _guard1736 = ev00__0state <= 6'd29;
wire _guard1737 = _guard1735 & _guard1736;
wire _guard1738 = _guard1734 | _guard1737;
wire _guard1739 = ev00__0state >= 6'd42;
wire _guard1740 = ev00__0state <= 6'd42;
wire _guard1741 = _guard1739 & _guard1740;
wire _guard1742 = _guard1738 | _guard1741;
wire _guard1743 = ev00__0state >= 6'd4;
wire _guard1744 = ev00__0state <= 6'd4;
wire _guard1745 = _guard1743 & _guard1744;
wire _guard1746 = _guard1742 | _guard1745;
wire _guard1747 = ev00__0state >= 6'd17;
wire _guard1748 = ev00__0state <= 6'd17;
wire _guard1749 = _guard1747 & _guard1748;
wire _guard1750 = _guard1746 | _guard1749;
wire _guard1751 = ev00__0state >= 6'd30;
wire _guard1752 = ev00__0state <= 6'd30;
wire _guard1753 = _guard1751 & _guard1752;
wire _guard1754 = _guard1750 | _guard1753;
wire _guard1755 = ev00__0state >= 6'd43;
wire _guard1756 = ev00__0state <= 6'd43;
wire _guard1757 = _guard1755 & _guard1756;
wire _guard1758 = _guard1754 | _guard1757;
wire _guard1759 = ev00__0state >= 6'd5;
wire _guard1760 = ev00__0state <= 6'd5;
wire _guard1761 = _guard1759 & _guard1760;
wire _guard1762 = _guard1758 | _guard1761;
wire _guard1763 = ev00__0state >= 6'd18;
wire _guard1764 = ev00__0state <= 6'd18;
wire _guard1765 = _guard1763 & _guard1764;
wire _guard1766 = _guard1762 | _guard1765;
wire _guard1767 = ev00__0state >= 6'd31;
wire _guard1768 = ev00__0state <= 6'd31;
wire _guard1769 = _guard1767 & _guard1768;
wire _guard1770 = _guard1766 | _guard1769;
wire _guard1771 = ev00__0state >= 6'd44;
wire _guard1772 = ev00__0state <= 6'd44;
wire _guard1773 = _guard1771 & _guard1772;
wire _guard1774 = _guard1770 | _guard1773;
wire _guard1775 = ev00__0state >= 6'd6;
wire _guard1776 = ev00__0state <= 6'd6;
wire _guard1777 = _guard1775 & _guard1776;
wire _guard1778 = _guard1774 | _guard1777;
wire _guard1779 = ev00__0state >= 6'd19;
wire _guard1780 = ev00__0state <= 6'd19;
wire _guard1781 = _guard1779 & _guard1780;
wire _guard1782 = _guard1778 | _guard1781;
wire _guard1783 = ev00__0state >= 6'd32;
wire _guard1784 = ev00__0state <= 6'd32;
wire _guard1785 = _guard1783 & _guard1784;
wire _guard1786 = _guard1782 | _guard1785;
wire _guard1787 = ev00__0state >= 6'd45;
wire _guard1788 = ev00__0state <= 6'd45;
wire _guard1789 = _guard1787 & _guard1788;
wire _guard1790 = _guard1786 | _guard1789;
wire _guard1791 = ev00__0state >= 6'd7;
wire _guard1792 = ev00__0state <= 6'd7;
wire _guard1793 = _guard1791 & _guard1792;
wire _guard1794 = _guard1790 | _guard1793;
wire _guard1795 = ev00__0state >= 6'd20;
wire _guard1796 = ev00__0state <= 6'd20;
wire _guard1797 = _guard1795 & _guard1796;
wire _guard1798 = _guard1794 | _guard1797;
wire _guard1799 = ev00__0state >= 6'd33;
wire _guard1800 = ev00__0state <= 6'd33;
wire _guard1801 = _guard1799 & _guard1800;
wire _guard1802 = _guard1798 | _guard1801;
wire _guard1803 = ev00__0state >= 6'd46;
wire _guard1804 = ev00__0state <= 6'd46;
wire _guard1805 = _guard1803 & _guard1804;
wire _guard1806 = _guard1802 | _guard1805;
wire _guard1807 = ev00__0state >= 6'd2;
wire _guard1808 = ev00__0state <= 6'd2;
wire _guard1809 = _guard1807 & _guard1808;
wire _guard1810 = ev00__0state >= 6'd41;
wire _guard1811 = ev00__0state <= 6'd41;
wire _guard1812 = _guard1810 & _guard1811;
wire _guard1813 = ev00__0state >= 6'd31;
wire _guard1814 = ev00__0state <= 6'd31;
wire _guard1815 = _guard1813 & _guard1814;
wire _guard1816 = ev00__0state >= 6'd43;
wire _guard1817 = ev00__0state <= 6'd43;
wire _guard1818 = _guard1816 & _guard1817;
wire _guard1819 = ev00__0state >= 6'd27;
wire _guard1820 = ev00__0state <= 6'd27;
wire _guard1821 = _guard1819 & _guard1820;
wire _guard1822 = ev00__0state >= 6'd3;
wire _guard1823 = ev00__0state <= 6'd3;
wire _guard1824 = _guard1822 & _guard1823;
wire _guard1825 = ev00__0state >= 6'd33;
wire _guard1826 = ev00__0state <= 6'd33;
wire _guard1827 = _guard1825 & _guard1826;
wire _guard1828 = ev00__0state >= 6'd14;
wire _guard1829 = ev00__0state <= 6'd14;
wire _guard1830 = _guard1828 & _guard1829;
wire _guard1831 = ev00__0state >= 6'd32;
wire _guard1832 = ev00__0state <= 6'd32;
wire _guard1833 = _guard1831 & _guard1832;
wire _guard1834 = ev00__0state >= 6'd5;
wire _guard1835 = ev00__0state <= 6'd5;
wire _guard1836 = _guard1834 & _guard1835;
wire _guard1837 = ev00__0state >= 6'd45;
wire _guard1838 = ev00__0state <= 6'd45;
wire _guard1839 = _guard1837 & _guard1838;
wire _guard1840 = ev00__0state >= 6'd40;
wire _guard1841 = ev00__0state <= 6'd40;
wire _guard1842 = _guard1840 & _guard1841;
wire _guard1843 = ev00__0state >= 6'd28;
wire _guard1844 = ev00__0state <= 6'd28;
wire _guard1845 = _guard1843 & _guard1844;
wire _guard1846 = ev00__0state >= 6'd17;
wire _guard1847 = ev00__0state <= 6'd17;
wire _guard1848 = _guard1846 & _guard1847;
wire _guard1849 = ev00__0state >= 6'd19;
wire _guard1850 = ev00__0state <= 6'd19;
wire _guard1851 = _guard1849 & _guard1850;
wire _guard1852 = ev00__0state >= 6'd15;
wire _guard1853 = ev00__0state <= 6'd15;
wire _guard1854 = _guard1852 & _guard1853;
wire _guard1855 = ev00__0state >= 6'd4;
wire _guard1856 = ev00__0state <= 6'd4;
wire _guard1857 = _guard1855 & _guard1856;
wire _guard1858 = ev00__0state >= 6'd46;
wire _guard1859 = ev00__0state <= 6'd46;
wire _guard1860 = _guard1858 & _guard1859;
wire _guard1861 = ev00__0state >= 6'd1;
wire _guard1862 = ev00__0state <= 6'd1;
wire _guard1863 = _guard1861 & _guard1862;
wire _guard1864 = ev00__0state >= 6'd16;
wire _guard1865 = ev00__0state <= 6'd16;
wire _guard1866 = _guard1864 & _guard1865;
wire _guard1867 = ev00__0state >= 6'd20;
wire _guard1868 = ev00__0state <= 6'd20;
wire _guard1869 = _guard1867 & _guard1868;
wire _guard1870 = ev00__0state >= 6'd7;
wire _guard1871 = ev00__0state <= 6'd7;
wire _guard1872 = _guard1870 & _guard1871;
wire _guard1873 = ev00__0state >= 6'd42;
wire _guard1874 = ev00__0state <= 6'd42;
wire _guard1875 = _guard1873 & _guard1874;
wire _guard1876 = ev00__0state >= 6'd29;
wire _guard1877 = ev00__0state <= 6'd29;
wire _guard1878 = _guard1876 & _guard1877;
wire _guard1879 = ev00__0state >= 6'd44;
wire _guard1880 = ev00__0state <= 6'd44;
wire _guard1881 = _guard1879 & _guard1880;
wire _guard1882 = ev00__0state >= 6'd6;
wire _guard1883 = ev00__0state <= 6'd6;
wire _guard1884 = _guard1882 & _guard1883;
wire _guard1885 = ev00__0state >= 6'd13;
wire _guard1886 = ev00__0state <= 6'd13;
wire _guard1887 = _guard1885 & _guard1886;
wire _guard1888 = ev00__0state >= 6'd26;
wire _guard1889 = ev00__0state <= 6'd26;
wire _guard1890 = _guard1888 & _guard1889;
wire _guard1891 = ev00__0state >= 6'd39;
wire _guard1892 = ev00__0state <= 6'd39;
wire _guard1893 = _guard1891 & _guard1892;
wire _guard1894 = ev00__0state >= 6'd30;
wire _guard1895 = ev00__0state <= 6'd30;
wire _guard1896 = _guard1894 & _guard1895;
wire _guard1897 = ev00__0_0;
wire _guard1898 = ev00__0state >= 6'd1;
wire _guard1899 = ev00__0state <= 6'd0;
wire _guard1900 = _guard1898 & _guard1899;
wire _guard1901 = _guard1897 | _guard1900;
wire _guard1902 = ev00__0state >= 6'd18;
wire _guard1903 = ev00__0state <= 6'd18;
wire _guard1904 = _guard1902 & _guard1903;
wire _guard1905 = ev00__0state >= 6'd2;
wire _guard1906 = ev00__0state <= 6'd2;
wire _guard1907 = _guard1905 & _guard1906;
wire _guard1908 = ev00__0state >= 6'd41;
wire _guard1909 = ev00__0state <= 6'd41;
wire _guard1910 = _guard1908 & _guard1909;
wire _guard1911 = ev00__0state >= 6'd31;
wire _guard1912 = ev00__0state <= 6'd31;
wire _guard1913 = _guard1911 & _guard1912;
wire _guard1914 = ev00__0state >= 6'd43;
wire _guard1915 = ev00__0state <= 6'd43;
wire _guard1916 = _guard1914 & _guard1915;
wire _guard1917 = ev00__0state >= 6'd27;
wire _guard1918 = ev00__0state <= 6'd27;
wire _guard1919 = _guard1917 & _guard1918;
wire _guard1920 = ev00__0state >= 6'd3;
wire _guard1921 = ev00__0state <= 6'd3;
wire _guard1922 = _guard1920 & _guard1921;
wire _guard1923 = ev00__0state >= 6'd33;
wire _guard1924 = ev00__0state <= 6'd33;
wire _guard1925 = _guard1923 & _guard1924;
wire _guard1926 = ev00__0state >= 6'd14;
wire _guard1927 = ev00__0state <= 6'd14;
wire _guard1928 = _guard1926 & _guard1927;
wire _guard1929 = ev00__0state >= 6'd32;
wire _guard1930 = ev00__0state <= 6'd32;
wire _guard1931 = _guard1929 & _guard1930;
wire _guard1932 = ev00__0state >= 6'd5;
wire _guard1933 = ev00__0state <= 6'd5;
wire _guard1934 = _guard1932 & _guard1933;
wire _guard1935 = ev00__0state >= 6'd45;
wire _guard1936 = ev00__0state <= 6'd45;
wire _guard1937 = _guard1935 & _guard1936;
wire _guard1938 = ev00__0state >= 6'd40;
wire _guard1939 = ev00__0state <= 6'd40;
wire _guard1940 = _guard1938 & _guard1939;
wire _guard1941 = ev00__0state >= 6'd28;
wire _guard1942 = ev00__0state <= 6'd28;
wire _guard1943 = _guard1941 & _guard1942;
wire _guard1944 = ev00__0state >= 6'd17;
wire _guard1945 = ev00__0state <= 6'd17;
wire _guard1946 = _guard1944 & _guard1945;
wire _guard1947 = ev00__0state >= 6'd19;
wire _guard1948 = ev00__0state <= 6'd19;
wire _guard1949 = _guard1947 & _guard1948;
wire _guard1950 = ev00__0state >= 6'd15;
wire _guard1951 = ev00__0state <= 6'd15;
wire _guard1952 = _guard1950 & _guard1951;
wire _guard1953 = ev00__0state >= 6'd4;
wire _guard1954 = ev00__0state <= 6'd4;
wire _guard1955 = _guard1953 & _guard1954;
wire _guard1956 = ev00__0state >= 6'd46;
wire _guard1957 = ev00__0state <= 6'd46;
wire _guard1958 = _guard1956 & _guard1957;
wire _guard1959 = ev00__0state >= 6'd1;
wire _guard1960 = ev00__0state <= 6'd1;
wire _guard1961 = _guard1959 & _guard1960;
wire _guard1962 = ev00__0state >= 6'd16;
wire _guard1963 = ev00__0state <= 6'd16;
wire _guard1964 = _guard1962 & _guard1963;
wire _guard1965 = ev00__0state >= 6'd20;
wire _guard1966 = ev00__0state <= 6'd20;
wire _guard1967 = _guard1965 & _guard1966;
wire _guard1968 = ev00__0state >= 6'd7;
wire _guard1969 = ev00__0state <= 6'd7;
wire _guard1970 = _guard1968 & _guard1969;
wire _guard1971 = ev00__0state >= 6'd42;
wire _guard1972 = ev00__0state <= 6'd42;
wire _guard1973 = _guard1971 & _guard1972;
wire _guard1974 = ev00__0state >= 6'd29;
wire _guard1975 = ev00__0state <= 6'd29;
wire _guard1976 = _guard1974 & _guard1975;
wire _guard1977 = ev00__0state >= 6'd44;
wire _guard1978 = ev00__0state <= 6'd44;
wire _guard1979 = _guard1977 & _guard1978;
wire _guard1980 = ev00__0state >= 6'd6;
wire _guard1981 = ev00__0state <= 6'd6;
wire _guard1982 = _guard1980 & _guard1981;
wire _guard1983 = ev00__0state >= 6'd13;
wire _guard1984 = ev00__0state <= 6'd13;
wire _guard1985 = _guard1983 & _guard1984;
wire _guard1986 = ev00__0state >= 6'd26;
wire _guard1987 = ev00__0state <= 6'd26;
wire _guard1988 = _guard1986 & _guard1987;
wire _guard1989 = ev00__0state >= 6'd39;
wire _guard1990 = ev00__0state <= 6'd39;
wire _guard1991 = _guard1989 & _guard1990;
wire _guard1992 = ev00__0state >= 6'd30;
wire _guard1993 = ev00__0state <= 6'd30;
wire _guard1994 = _guard1992 & _guard1993;
wire _guard1995 = ev00__0_0;
wire _guard1996 = ev00__0state >= 6'd1;
wire _guard1997 = ev00__0state <= 6'd0;
wire _guard1998 = _guard1996 & _guard1997;
wire _guard1999 = _guard1995 | _guard1998;
wire _guard2000 = ev00__0state >= 6'd18;
wire _guard2001 = ev00__0state <= 6'd18;
wire _guard2002 = _guard2000 & _guard2001;
wire _guard2003 = ev00__0state >= 6'd2;
wire _guard2004 = ev00__0state <= 6'd2;
wire _guard2005 = _guard2003 & _guard2004;
wire _guard2006 = ev00__0state >= 6'd41;
wire _guard2007 = ev00__0state <= 6'd41;
wire _guard2008 = _guard2006 & _guard2007;
wire _guard2009 = ev00__0state >= 6'd31;
wire _guard2010 = ev00__0state <= 6'd31;
wire _guard2011 = _guard2009 & _guard2010;
wire _guard2012 = ev00__0state >= 6'd43;
wire _guard2013 = ev00__0state <= 6'd43;
wire _guard2014 = _guard2012 & _guard2013;
wire _guard2015 = ev00__0state >= 6'd27;
wire _guard2016 = ev00__0state <= 6'd27;
wire _guard2017 = _guard2015 & _guard2016;
wire _guard2018 = ev00__0state >= 6'd3;
wire _guard2019 = ev00__0state <= 6'd3;
wire _guard2020 = _guard2018 & _guard2019;
wire _guard2021 = ev00__0state >= 6'd33;
wire _guard2022 = ev00__0state <= 6'd33;
wire _guard2023 = _guard2021 & _guard2022;
wire _guard2024 = ev00__0state >= 6'd14;
wire _guard2025 = ev00__0state <= 6'd14;
wire _guard2026 = _guard2024 & _guard2025;
wire _guard2027 = ev00__0state >= 6'd32;
wire _guard2028 = ev00__0state <= 6'd32;
wire _guard2029 = _guard2027 & _guard2028;
wire _guard2030 = ev00__0state >= 6'd5;
wire _guard2031 = ev00__0state <= 6'd5;
wire _guard2032 = _guard2030 & _guard2031;
wire _guard2033 = ev00__0state >= 6'd45;
wire _guard2034 = ev00__0state <= 6'd45;
wire _guard2035 = _guard2033 & _guard2034;
wire _guard2036 = ev00__0state >= 6'd40;
wire _guard2037 = ev00__0state <= 6'd40;
wire _guard2038 = _guard2036 & _guard2037;
wire _guard2039 = ev00__0state >= 6'd28;
wire _guard2040 = ev00__0state <= 6'd28;
wire _guard2041 = _guard2039 & _guard2040;
wire _guard2042 = ev00__0state >= 6'd17;
wire _guard2043 = ev00__0state <= 6'd17;
wire _guard2044 = _guard2042 & _guard2043;
wire _guard2045 = ev00__0state >= 6'd19;
wire _guard2046 = ev00__0state <= 6'd19;
wire _guard2047 = _guard2045 & _guard2046;
wire _guard2048 = ev00__0state >= 6'd15;
wire _guard2049 = ev00__0state <= 6'd15;
wire _guard2050 = _guard2048 & _guard2049;
wire _guard2051 = ev00__0state >= 6'd4;
wire _guard2052 = ev00__0state <= 6'd4;
wire _guard2053 = _guard2051 & _guard2052;
wire _guard2054 = ev00__0state >= 6'd46;
wire _guard2055 = ev00__0state <= 6'd46;
wire _guard2056 = _guard2054 & _guard2055;
wire _guard2057 = ev00__0state >= 6'd1;
wire _guard2058 = ev00__0state <= 6'd1;
wire _guard2059 = _guard2057 & _guard2058;
wire _guard2060 = ev00__0state >= 6'd16;
wire _guard2061 = ev00__0state <= 6'd16;
wire _guard2062 = _guard2060 & _guard2061;
wire _guard2063 = ev00__0state >= 6'd20;
wire _guard2064 = ev00__0state <= 6'd20;
wire _guard2065 = _guard2063 & _guard2064;
wire _guard2066 = ev00__0state >= 6'd7;
wire _guard2067 = ev00__0state <= 6'd7;
wire _guard2068 = _guard2066 & _guard2067;
wire _guard2069 = ev00__0state >= 6'd42;
wire _guard2070 = ev00__0state <= 6'd42;
wire _guard2071 = _guard2069 & _guard2070;
wire _guard2072 = ev00__0state >= 6'd29;
wire _guard2073 = ev00__0state <= 6'd29;
wire _guard2074 = _guard2072 & _guard2073;
wire _guard2075 = ev00__0state >= 6'd44;
wire _guard2076 = ev00__0state <= 6'd44;
wire _guard2077 = _guard2075 & _guard2076;
wire _guard2078 = ev00__0state >= 6'd6;
wire _guard2079 = ev00__0state <= 6'd6;
wire _guard2080 = _guard2078 & _guard2079;
wire _guard2081 = ev00__0state >= 6'd13;
wire _guard2082 = ev00__0state <= 6'd13;
wire _guard2083 = _guard2081 & _guard2082;
wire _guard2084 = ev00__0state >= 6'd26;
wire _guard2085 = ev00__0state <= 6'd26;
wire _guard2086 = _guard2084 & _guard2085;
wire _guard2087 = ev00__0state >= 6'd39;
wire _guard2088 = ev00__0state <= 6'd39;
wire _guard2089 = _guard2087 & _guard2088;
wire _guard2090 = ev00__0state >= 6'd30;
wire _guard2091 = ev00__0state <= 6'd30;
wire _guard2092 = _guard2090 & _guard2091;
wire _guard2093 = ev00__0_0;
wire _guard2094 = ev00__0state >= 6'd1;
wire _guard2095 = ev00__0state <= 6'd0;
wire _guard2096 = _guard2094 & _guard2095;
wire _guard2097 = _guard2093 | _guard2096;
wire _guard2098 = ev00__0state >= 6'd18;
wire _guard2099 = ev00__0state <= 6'd18;
wire _guard2100 = _guard2098 & _guard2099;
wire _guard2101 = ev00__0state >= 6'd2;
wire _guard2102 = ev00__0state <= 6'd2;
wire _guard2103 = _guard2101 & _guard2102;
wire _guard2104 = ev00__0state >= 6'd41;
wire _guard2105 = ev00__0state <= 6'd41;
wire _guard2106 = _guard2104 & _guard2105;
wire _guard2107 = ev00__0state >= 6'd31;
wire _guard2108 = ev00__0state <= 6'd31;
wire _guard2109 = _guard2107 & _guard2108;
wire _guard2110 = ev00__0state >= 6'd43;
wire _guard2111 = ev00__0state <= 6'd43;
wire _guard2112 = _guard2110 & _guard2111;
wire _guard2113 = ev00__0state >= 6'd27;
wire _guard2114 = ev00__0state <= 6'd27;
wire _guard2115 = _guard2113 & _guard2114;
wire _guard2116 = ev00__0state >= 6'd3;
wire _guard2117 = ev00__0state <= 6'd3;
wire _guard2118 = _guard2116 & _guard2117;
wire _guard2119 = ev00__0state >= 6'd33;
wire _guard2120 = ev00__0state <= 6'd33;
wire _guard2121 = _guard2119 & _guard2120;
wire _guard2122 = ev00__0state >= 6'd14;
wire _guard2123 = ev00__0state <= 6'd14;
wire _guard2124 = _guard2122 & _guard2123;
wire _guard2125 = ev00__0state >= 6'd32;
wire _guard2126 = ev00__0state <= 6'd32;
wire _guard2127 = _guard2125 & _guard2126;
wire _guard2128 = ev00__0state >= 6'd5;
wire _guard2129 = ev00__0state <= 6'd5;
wire _guard2130 = _guard2128 & _guard2129;
wire _guard2131 = ev00__0state >= 6'd45;
wire _guard2132 = ev00__0state <= 6'd45;
wire _guard2133 = _guard2131 & _guard2132;
wire _guard2134 = ev00__0state >= 6'd40;
wire _guard2135 = ev00__0state <= 6'd40;
wire _guard2136 = _guard2134 & _guard2135;
wire _guard2137 = ev00__0state >= 6'd28;
wire _guard2138 = ev00__0state <= 6'd28;
wire _guard2139 = _guard2137 & _guard2138;
wire _guard2140 = ev00__0state >= 6'd17;
wire _guard2141 = ev00__0state <= 6'd17;
wire _guard2142 = _guard2140 & _guard2141;
wire _guard2143 = ev00__0state >= 6'd19;
wire _guard2144 = ev00__0state <= 6'd19;
wire _guard2145 = _guard2143 & _guard2144;
wire _guard2146 = ev00__0state >= 6'd15;
wire _guard2147 = ev00__0state <= 6'd15;
wire _guard2148 = _guard2146 & _guard2147;
wire _guard2149 = ev00__0state >= 6'd4;
wire _guard2150 = ev00__0state <= 6'd4;
wire _guard2151 = _guard2149 & _guard2150;
wire _guard2152 = ev00__0state >= 6'd46;
wire _guard2153 = ev00__0state <= 6'd46;
wire _guard2154 = _guard2152 & _guard2153;
wire _guard2155 = ev00__0state >= 6'd1;
wire _guard2156 = ev00__0state <= 6'd1;
wire _guard2157 = _guard2155 & _guard2156;
wire _guard2158 = ev00__0state >= 6'd16;
wire _guard2159 = ev00__0state <= 6'd16;
wire _guard2160 = _guard2158 & _guard2159;
wire _guard2161 = ev00__0state >= 6'd20;
wire _guard2162 = ev00__0state <= 6'd20;
wire _guard2163 = _guard2161 & _guard2162;
wire _guard2164 = ev00__0state >= 6'd7;
wire _guard2165 = ev00__0state <= 6'd7;
wire _guard2166 = _guard2164 & _guard2165;
wire _guard2167 = ev00__0state >= 6'd42;
wire _guard2168 = ev00__0state <= 6'd42;
wire _guard2169 = _guard2167 & _guard2168;
wire _guard2170 = ev00__0state >= 6'd29;
wire _guard2171 = ev00__0state <= 6'd29;
wire _guard2172 = _guard2170 & _guard2171;
wire _guard2173 = ev00__0state >= 6'd44;
wire _guard2174 = ev00__0state <= 6'd44;
wire _guard2175 = _guard2173 & _guard2174;
wire _guard2176 = ev00__0state >= 6'd6;
wire _guard2177 = ev00__0state <= 6'd6;
wire _guard2178 = _guard2176 & _guard2177;
wire _guard2179 = ev00__0state >= 6'd13;
wire _guard2180 = ev00__0state <= 6'd13;
wire _guard2181 = _guard2179 & _guard2180;
wire _guard2182 = ev00__0state >= 6'd26;
wire _guard2183 = ev00__0state <= 6'd26;
wire _guard2184 = _guard2182 & _guard2183;
wire _guard2185 = ev00__0state >= 6'd39;
wire _guard2186 = ev00__0state <= 6'd39;
wire _guard2187 = _guard2185 & _guard2186;
wire _guard2188 = ev00__0state >= 6'd30;
wire _guard2189 = ev00__0state <= 6'd30;
wire _guard2190 = _guard2188 & _guard2189;
wire _guard2191 = ev00__0_0;
wire _guard2192 = ev00__0state >= 6'd1;
wire _guard2193 = ev00__0state <= 6'd0;
wire _guard2194 = _guard2192 & _guard2193;
wire _guard2195 = _guard2191 | _guard2194;
wire _guard2196 = ev00__0state >= 6'd18;
wire _guard2197 = ev00__0state <= 6'd18;
wire _guard2198 = _guard2196 & _guard2197;
wire _guard2199 = ev00__0_0;
wire _guard2200 = ev00__0state >= 6'd1;
wire _guard2201 = ev00__0state <= 6'd0;
wire _guard2202 = _guard2200 & _guard2201;
wire _guard2203 = _guard2199 | _guard2202;
wire _guard2204 = ev00__0state >= 6'd5;
wire _guard2205 = ev00__0state <= 6'd5;
wire _guard2206 = _guard2204 & _guard2205;
wire _guard2207 = ev00__0state >= 6'd1;
wire _guard2208 = ev00__0state <= 6'd1;
wire _guard2209 = _guard2207 & _guard2208;
wire _guard2210 = ev00__0state >= 6'd2;
wire _guard2211 = ev00__0state <= 6'd2;
wire _guard2212 = _guard2210 & _guard2211;
wire _guard2213 = ev00__0state >= 6'd3;
wire _guard2214 = ev00__0state <= 6'd3;
wire _guard2215 = _guard2213 & _guard2214;
wire _guard2216 = ev00__0state >= 6'd6;
wire _guard2217 = ev00__0state <= 6'd6;
wire _guard2218 = _guard2216 & _guard2217;
wire _guard2219 = ev00__0state >= 6'd4;
wire _guard2220 = ev00__0state <= 6'd4;
wire _guard2221 = _guard2219 & _guard2220;
wire _guard2222 = ev00__0state >= 6'd7;
wire _guard2223 = ev00__0state <= 6'd7;
wire _guard2224 = _guard2222 & _guard2223;
wire _guard2225 = ev00__0state >= 6'd39;
wire _guard2226 = ev00__0state <= 6'd39;
wire _guard2227 = _guard2225 & _guard2226;
wire _guard2228 = ev00__0state >= 6'd44;
wire _guard2229 = ev00__0state <= 6'd44;
wire _guard2230 = _guard2228 & _guard2229;
wire _guard2231 = ev00__0state >= 6'd40;
wire _guard2232 = ev00__0state <= 6'd40;
wire _guard2233 = _guard2231 & _guard2232;
wire _guard2234 = ev00__0state >= 6'd41;
wire _guard2235 = ev00__0state <= 6'd41;
wire _guard2236 = _guard2234 & _guard2235;
wire _guard2237 = ev00__0state >= 6'd42;
wire _guard2238 = ev00__0state <= 6'd42;
wire _guard2239 = _guard2237 & _guard2238;
wire _guard2240 = ev00__0state >= 6'd45;
wire _guard2241 = ev00__0state <= 6'd45;
wire _guard2242 = _guard2240 & _guard2241;
wire _guard2243 = ev00__0state >= 6'd43;
wire _guard2244 = ev00__0state <= 6'd43;
wire _guard2245 = _guard2243 & _guard2244;
wire _guard2246 = ev00__0state >= 6'd46;
wire _guard2247 = ev00__0state <= 6'd46;
wire _guard2248 = _guard2246 & _guard2247;
wire _guard2249 = ev00__0state >= 6'd26;
wire _guard2250 = ev00__0state <= 6'd26;
wire _guard2251 = _guard2249 & _guard2250;
wire _guard2252 = ev00__0state >= 6'd31;
wire _guard2253 = ev00__0state <= 6'd31;
wire _guard2254 = _guard2252 & _guard2253;
wire _guard2255 = ev00__0state >= 6'd27;
wire _guard2256 = ev00__0state <= 6'd27;
wire _guard2257 = _guard2255 & _guard2256;
wire _guard2258 = ev00__0state >= 6'd28;
wire _guard2259 = ev00__0state <= 6'd28;
wire _guard2260 = _guard2258 & _guard2259;
wire _guard2261 = ev00__0state >= 6'd29;
wire _guard2262 = ev00__0state <= 6'd29;
wire _guard2263 = _guard2261 & _guard2262;
wire _guard2264 = ev00__0state >= 6'd32;
wire _guard2265 = ev00__0state <= 6'd32;
wire _guard2266 = _guard2264 & _guard2265;
wire _guard2267 = ev00__0state >= 6'd30;
wire _guard2268 = ev00__0state <= 6'd30;
wire _guard2269 = _guard2267 & _guard2268;
wire _guard2270 = ev00__0state >= 6'd33;
wire _guard2271 = ev00__0state <= 6'd33;
wire _guard2272 = _guard2270 & _guard2271;
wire _guard2273 = ev00__0state >= 6'd13;
wire _guard2274 = ev00__0state <= 6'd13;
wire _guard2275 = _guard2273 & _guard2274;
wire _guard2276 = ev00__0state >= 6'd18;
wire _guard2277 = ev00__0state <= 6'd18;
wire _guard2278 = _guard2276 & _guard2277;
wire _guard2279 = ev00__0state >= 6'd14;
wire _guard2280 = ev00__0state <= 6'd14;
wire _guard2281 = _guard2279 & _guard2280;
wire _guard2282 = ev00__0state >= 6'd15;
wire _guard2283 = ev00__0state <= 6'd15;
wire _guard2284 = _guard2282 & _guard2283;
wire _guard2285 = ev00__0state >= 6'd16;
wire _guard2286 = ev00__0state <= 6'd16;
wire _guard2287 = _guard2285 & _guard2286;
wire _guard2288 = ev00__0state >= 6'd19;
wire _guard2289 = ev00__0state <= 6'd19;
wire _guard2290 = _guard2288 & _guard2289;
wire _guard2291 = ev00__0state >= 6'd17;
wire _guard2292 = ev00__0state <= 6'd17;
wire _guard2293 = _guard2291 & _guard2292;
wire _guard2294 = ev00__0state >= 6'd20;
wire _guard2295 = ev00__0state <= 6'd20;
wire _guard2296 = _guard2294 & _guard2295;
wire _guard2297 = ev00__0_0;
wire _guard2298 = ev00__0state >= 6'd1;
wire _guard2299 = ev00__0state <= 6'd51;
wire _guard2300 = _guard2298 & _guard2299;
wire _guard2301 = _guard2297 | _guard2300;
wire _guard2302 = ev00__0_0;
wire _guard2303 = ev00__0state >= 6'd1;
wire _guard2304 = ev00__0state <= 6'd51;
wire _guard2305 = _guard2303 & _guard2304;
wire _guard2306 = _guard2302 | _guard2305;
wire _guard2307 = ev00__0_0;
wire _guard2308 = ev00__0state >= 6'd1;
wire _guard2309 = ev00__0state <= 6'd51;
wire _guard2310 = _guard2308 & _guard2309;
wire _guard2311 = _guard2307 | _guard2310;
wire _guard2312 = ev00__0_0;
wire _guard2313 = ev00__0state >= 6'd1;
wire _guard2314 = ev00__0state <= 6'd51;
wire _guard2315 = _guard2313 & _guard2314;
wire _guard2316 = _guard2312 | _guard2315;
wire _guard2317 = ev00__0_0;
wire _guard2318 = ev00__0state >= 6'd1;
wire _guard2319 = ev00__0state <= 6'd51;
wire _guard2320 = _guard2318 & _guard2319;
wire _guard2321 = _guard2317 | _guard2320;
wire _guard2322 = ev00__0_0;
wire _guard2323 = ev00__0state >= 6'd1;
wire _guard2324 = ev00__0state <= 6'd51;
wire _guard2325 = _guard2323 & _guard2324;
wire _guard2326 = _guard2322 | _guard2325;
wire _guard2327 = ev00__0_0;
wire _guard2328 = ev00__0state >= 6'd1;
wire _guard2329 = ev00__0state <= 6'd51;
wire _guard2330 = _guard2328 & _guard2329;
wire _guard2331 = _guard2327 | _guard2330;
wire _guard2332 = ev00__0_0;
wire _guard2333 = ev00__0state >= 6'd1;
wire _guard2334 = ev00__0state <= 6'd51;
wire _guard2335 = _guard2333 & _guard2334;
wire _guard2336 = _guard2332 | _guard2335;
wire _guard2337 = ev00__0_0;
wire _guard2338 = ev00__0state >= 6'd1;
wire _guard2339 = ev00__0state <= 6'd51;
wire _guard2340 = _guard2338 & _guard2339;
wire _guard2341 = _guard2337 | _guard2340;
wire _guard2342 = ev00__0_0;
wire _guard2343 = ev00__0state >= 6'd1;
wire _guard2344 = ev00__0state <= 6'd51;
wire _guard2345 = _guard2343 & _guard2344;
wire _guard2346 = _guard2342 | _guard2345;
wire _guard2347 = ev00__0_0;
wire _guard2348 = ev00__0state >= 6'd1;
wire _guard2349 = ev00__0state <= 6'd51;
wire _guard2350 = _guard2348 & _guard2349;
wire _guard2351 = _guard2347 | _guard2350;
wire _guard2352 = ev00__0_0;
wire _guard2353 = ev00__0state >= 6'd1;
wire _guard2354 = ev00__0state <= 6'd51;
wire _guard2355 = _guard2353 & _guard2354;
wire _guard2356 = _guard2352 | _guard2355;
wire _guard2357 = ev00__0_0;
wire _guard2358 = ev00__0state >= 6'd1;
wire _guard2359 = ev00__0state <= 6'd51;
wire _guard2360 = _guard2358 & _guard2359;
wire _guard2361 = _guard2357 | _guard2360;
wire _guard2362 = ev00__0_0;
wire _guard2363 = ev00__0state >= 6'd1;
wire _guard2364 = ev00__0state <= 6'd51;
wire _guard2365 = _guard2363 & _guard2364;
wire _guard2366 = _guard2362 | _guard2365;
wire _guard2367 = ev00__0_0;
wire _guard2368 = ev00__0state >= 6'd1;
wire _guard2369 = ev00__0state <= 6'd51;
wire _guard2370 = _guard2368 & _guard2369;
wire _guard2371 = _guard2367 | _guard2370;
wire _guard2372 = ev00__0_0;
wire _guard2373 = ev00__0state >= 6'd1;
wire _guard2374 = ev00__0state <= 6'd51;
wire _guard2375 = _guard2373 & _guard2374;
wire _guard2376 = _guard2372 | _guard2375;
wire _guard2377 = ev00__0state >= 6'd39;
wire _guard2378 = ev00__0state <= 6'd39;
wire _guard2379 = _guard2377 & _guard2378;
wire _guard2380 = ev00__0state >= 6'd39;
wire _guard2381 = ev00__0state <= 6'd39;
wire _guard2382 = _guard2380 & _guard2381;
wire _guard2383 = ev00__0state >= 6'd39;
wire _guard2384 = ev00__0state <= 6'd39;
wire _guard2385 = _guard2383 & _guard2384;
wire _guard2386 = ev00__0state >= 6'd39;
wire _guard2387 = ev00__0state <= 6'd39;
wire _guard2388 = _guard2386 & _guard2387;
wire _guard2389 = ev00__0state >= 6'd1;
wire _guard2390 = ev00__0state <= 6'd1;
wire _guard2391 = _guard2389 & _guard2390;
wire _guard2392 = ev00__0state >= 6'd12;
wire _guard2393 = ev00__0state <= 6'd12;
wire _guard2394 = _guard2392 & _guard2393;
wire _guard2395 = ev00__0state >= 6'd39;
wire _guard2396 = ev00__0state <= 6'd39;
wire _guard2397 = _guard2395 & _guard2396;
wire _guard2398 = ev00__0state >= 6'd39;
wire _guard2399 = ev00__0state <= 6'd39;
wire _guard2400 = _guard2398 & _guard2399;
wire _guard2401 = ev00__0state >= 6'd39;
wire _guard2402 = ev00__0state <= 6'd39;
wire _guard2403 = _guard2401 & _guard2402;
wire _guard2404 = ev00__0state >= 6'd39;
wire _guard2405 = ev00__0state <= 6'd39;
wire _guard2406 = _guard2404 & _guard2405;
wire _guard2407 = ev00__0state >= 6'd51;
wire _guard2408 = ev00__0state <= 6'd51;
wire _guard2409 = _guard2407 & _guard2408;
wire _guard2410 = ev00__0state >= 6'd16;
wire _guard2411 = ev00__0state <= 6'd16;
wire _guard2412 = _guard2410 & _guard2411;
wire _guard2413 = ev00__0state >= 6'd8;
wire _guard2414 = ev00__0state <= 6'd8;
wire _guard2415 = _guard2413 & _guard2414;
wire _guard2416 = ev00__0state >= 6'd8;
wire _guard2417 = ev00__0state <= 6'd8;
wire _guard2418 = _guard2416 & _guard2417;
wire _guard2419 = ev00__0state >= 6'd8;
wire _guard2420 = ev00__0state <= 6'd8;
wire _guard2421 = _guard2419 & _guard2420;
wire _guard2422 = ev00__0state >= 6'd8;
wire _guard2423 = ev00__0state <= 6'd8;
wire _guard2424 = _guard2422 & _guard2423;
wire _guard2425 = ev00__0state >= 6'd10;
wire _guard2426 = ev00__0state <= 6'd10;
wire _guard2427 = _guard2425 & _guard2426;
wire _guard2428 = ev00__0state >= 6'd10;
wire _guard2429 = ev00__0state <= 6'd10;
wire _guard2430 = _guard2428 & _guard2429;
wire _guard2431 = ev00__0state >= 6'd10;
wire _guard2432 = ev00__0state <= 6'd10;
wire _guard2433 = _guard2431 & _guard2432;
wire _guard2434 = ev00__0state >= 6'd10;
wire _guard2435 = ev00__0state <= 6'd10;
wire _guard2436 = _guard2434 & _guard2435;
wire _guard2437 = ev00__0state >= 6'd49;
wire _guard2438 = ev00__0state <= 6'd49;
wire _guard2439 = _guard2437 & _guard2438;
wire _guard2440 = ev00__0state >= 6'd49;
wire _guard2441 = ev00__0state <= 6'd49;
wire _guard2442 = _guard2440 & _guard2441;
wire _guard2443 = ev00__0state >= 6'd49;
wire _guard2444 = ev00__0state <= 6'd49;
wire _guard2445 = _guard2443 & _guard2444;
wire _guard2446 = ev00__0state >= 6'd49;
wire _guard2447 = ev00__0state <= 6'd49;
wire _guard2448 = _guard2446 & _guard2447;
wire _guard2449 = ev00__0_0;
wire _guard2450 = ev00__0state >= 6'd1;
wire _guard2451 = ev00__0state <= 6'd0;
wire _guard2452 = _guard2450 & _guard2451;
wire _guard2453 = _guard2449 | _guard2452;
wire _guard2454 = ev00__0_0;
wire _guard2455 = ev00__0state >= 6'd1;
wire _guard2456 = ev00__0state <= 6'd0;
wire _guard2457 = _guard2455 & _guard2456;
wire _guard2458 = _guard2454 | _guard2457;
wire _guard2459 = ev00__0_0;
wire _guard2460 = ev00__0state >= 6'd1;
wire _guard2461 = ev00__0state <= 6'd0;
wire _guard2462 = _guard2460 & _guard2461;
wire _guard2463 = _guard2459 | _guard2462;
wire _guard2464 = ev00__0_0;
wire _guard2465 = ev00__0state >= 6'd1;
wire _guard2466 = ev00__0state <= 6'd0;
wire _guard2467 = _guard2465 & _guard2466;
wire _guard2468 = _guard2464 | _guard2467;
wire _guard2469 = ev00__0state >= 6'd20;
wire _guard2470 = ev00__0state <= 6'd20;
wire _guard2471 = _guard2469 & _guard2470;
wire _guard2472 = ev00__0state >= 6'd24;
wire _guard2473 = ev00__0state <= 6'd24;
wire _guard2474 = _guard2472 & _guard2473;
wire _guard2475 = ev00__0state >= 6'd24;
wire _guard2476 = ev00__0state <= 6'd24;
wire _guard2477 = _guard2475 & _guard2476;
wire _guard2478 = ev00__0state >= 6'd24;
wire _guard2479 = ev00__0state <= 6'd24;
wire _guard2480 = _guard2478 & _guard2479;
wire _guard2481 = ev00__0state >= 6'd24;
wire _guard2482 = ev00__0state <= 6'd24;
wire _guard2483 = _guard2481 & _guard2482;
wire _guard2484 = ev00__0state >= 6'd39;
wire _guard2485 = ev00__0state <= 6'd39;
wire _guard2486 = _guard2484 & _guard2485;
wire _guard2487 = ev00__0state >= 6'd39;
wire _guard2488 = ev00__0state <= 6'd39;
wire _guard2489 = _guard2487 & _guard2488;
wire _guard2490 = ev00__0state >= 6'd39;
wire _guard2491 = ev00__0state <= 6'd39;
wire _guard2492 = _guard2490 & _guard2491;
wire _guard2493 = ev00__0state >= 6'd39;
wire _guard2494 = ev00__0state <= 6'd39;
wire _guard2495 = _guard2493 & _guard2494;
wire _guard2496 = ev00__0state >= 6'd13;
wire _guard2497 = ev00__0state <= 6'd13;
wire _guard2498 = _guard2496 & _guard2497;
wire _guard2499 = ev00__0state >= 6'd26;
wire _guard2500 = ev00__0state <= 6'd26;
wire _guard2501 = _guard2499 & _guard2500;
wire _guard2502 = ev00__0state >= 6'd26;
wire _guard2503 = ev00__0state <= 6'd26;
wire _guard2504 = _guard2502 & _guard2503;
wire _guard2505 = ev00__0state >= 6'd26;
wire _guard2506 = ev00__0state <= 6'd26;
wire _guard2507 = _guard2505 & _guard2506;
wire _guard2508 = ev00__0state >= 6'd26;
wire _guard2509 = ev00__0state <= 6'd26;
wire _guard2510 = _guard2508 & _guard2509;
wire _guard2511 = ev00__0state >= 6'd39;
wire _guard2512 = ev00__0state <= 6'd39;
wire _guard2513 = _guard2511 & _guard2512;
wire _guard2514 = ev00__0state >= 6'd39;
wire _guard2515 = ev00__0state <= 6'd39;
wire _guard2516 = _guard2514 & _guard2515;
wire _guard2517 = ev00__0state >= 6'd39;
wire _guard2518 = ev00__0state <= 6'd39;
wire _guard2519 = _guard2517 & _guard2518;
wire _guard2520 = ev00__0state >= 6'd39;
wire _guard2521 = ev00__0state <= 6'd39;
wire _guard2522 = _guard2520 & _guard2521;
wire _guard2523 = ev00__0state >= 6'd12;
wire _guard2524 = ev00__0state <= 6'd12;
wire _guard2525 = _guard2523 & _guard2524;
wire _guard2526 = ev00__0state >= 6'd13;
wire _guard2527 = ev00__0state <= 6'd13;
wire _guard2528 = _guard2526 & _guard2527;
wire _guard2529 = ev00__0state >= 6'd13;
wire _guard2530 = ev00__0state <= 6'd13;
wire _guard2531 = _guard2529 & _guard2530;
wire _guard2532 = ev00__0state >= 6'd13;
wire _guard2533 = ev00__0state <= 6'd13;
wire _guard2534 = _guard2532 & _guard2533;
wire _guard2535 = ev00__0state >= 6'd13;
wire _guard2536 = ev00__0state <= 6'd13;
wire _guard2537 = _guard2535 & _guard2536;
wire _guard2538 = ev00__0state >= 6'd48;
wire _guard2539 = ev00__0state <= 6'd48;
wire _guard2540 = _guard2538 & _guard2539;
wire _guard2541 = ev00__0state >= 6'd48;
wire _guard2542 = ev00__0state <= 6'd48;
wire _guard2543 = _guard2541 & _guard2542;
wire _guard2544 = ev00__0state >= 6'd48;
wire _guard2545 = ev00__0state <= 6'd48;
wire _guard2546 = _guard2544 & _guard2545;
wire _guard2547 = ev00__0state >= 6'd48;
wire _guard2548 = ev00__0state <= 6'd48;
wire _guard2549 = _guard2547 & _guard2548;
wire _guard2550 = ev00__0state >= 6'd7;
wire _guard2551 = ev00__0state <= 6'd7;
wire _guard2552 = _guard2550 & _guard2551;
wire _guard2553 = ev00__0state >= 6'd32;
wire _guard2554 = ev00__0state <= 6'd32;
wire _guard2555 = _guard2553 & _guard2554;
wire _guard2556 = ev00__0state >= 6'd32;
wire _guard2557 = ev00__0state <= 6'd32;
wire _guard2558 = _guard2556 & _guard2557;
wire _guard2559 = ev00__0state >= 6'd32;
wire _guard2560 = ev00__0state <= 6'd32;
wire _guard2561 = _guard2559 & _guard2560;
wire _guard2562 = ev00__0state >= 6'd32;
wire _guard2563 = ev00__0state <= 6'd32;
wire _guard2564 = _guard2562 & _guard2563;
wire _guard2565 = ev00__0state >= 6'd42;
wire _guard2566 = ev00__0state <= 6'd42;
wire _guard2567 = _guard2565 & _guard2566;
wire _guard2568 = ev00__0state >= 6'd34;
wire _guard2569 = ev00__0state <= 6'd34;
wire _guard2570 = _guard2568 & _guard2569;
wire _guard2571 = ev00__0state >= 6'd34;
wire _guard2572 = ev00__0state <= 6'd34;
wire _guard2573 = _guard2571 & _guard2572;
wire _guard2574 = ev00__0state >= 6'd34;
wire _guard2575 = ev00__0state <= 6'd34;
wire _guard2576 = _guard2574 & _guard2575;
wire _guard2577 = ev00__0state >= 6'd34;
wire _guard2578 = ev00__0state <= 6'd34;
wire _guard2579 = _guard2577 & _guard2578;
wire _guard2580 = ev00__0state >= 6'd12;
wire _guard2581 = ev00__0state <= 6'd12;
wire _guard2582 = _guard2580 & _guard2581;
wire _guard2583 = ev00__0state >= 6'd25;
wire _guard2584 = ev00__0state <= 6'd25;
wire _guard2585 = _guard2583 & _guard2584;
wire _guard2586 = ev00__0_0;
wire _guard2587 = ev00__0state >= 6'd1;
wire _guard2588 = ev00__0state <= 6'd0;
wire _guard2589 = _guard2587 & _guard2588;
wire _guard2590 = _guard2586 | _guard2589;
wire _guard2591 = ev00__0_0;
wire _guard2592 = ev00__0state >= 6'd1;
wire _guard2593 = ev00__0state <= 6'd0;
wire _guard2594 = _guard2592 & _guard2593;
wire _guard2595 = _guard2591 | _guard2594;
wire _guard2596 = ev00__0_0;
wire _guard2597 = ev00__0state >= 6'd1;
wire _guard2598 = ev00__0state <= 6'd0;
wire _guard2599 = _guard2597 & _guard2598;
wire _guard2600 = _guard2596 | _guard2599;
wire _guard2601 = ev00__0_0;
wire _guard2602 = ev00__0state >= 6'd1;
wire _guard2603 = ev00__0state <= 6'd0;
wire _guard2604 = _guard2602 & _guard2603;
wire _guard2605 = _guard2601 | _guard2604;
wire _guard2606 = ev00__0state >= 6'd6;
wire _guard2607 = ev00__0state <= 6'd6;
wire _guard2608 = _guard2606 & _guard2607;
wire _guard2609 = ev00__0state >= 6'd6;
wire _guard2610 = ev00__0state <= 6'd6;
wire _guard2611 = _guard2609 & _guard2610;
wire _guard2612 = ev00__0state >= 6'd6;
wire _guard2613 = ev00__0state <= 6'd6;
wire _guard2614 = _guard2612 & _guard2613;
wire _guard2615 = ev00__0state >= 6'd6;
wire _guard2616 = ev00__0state <= 6'd6;
wire _guard2617 = _guard2615 & _guard2616;
wire _guard2618 = ev00__0state >= 6'd12;
wire _guard2619 = ev00__0state <= 6'd12;
wire _guard2620 = _guard2618 & _guard2619;
wire _guard2621 = ev00__0state >= 6'd29;
wire _guard2622 = ev00__0state <= 6'd29;
wire _guard2623 = _guard2621 & _guard2622;
wire _guard2624 = ev00__0state >= 6'd21;
wire _guard2625 = ev00__0state <= 6'd21;
wire _guard2626 = _guard2624 & _guard2625;
wire _guard2627 = ev00__0state >= 6'd21;
wire _guard2628 = ev00__0state <= 6'd21;
wire _guard2629 = _guard2627 & _guard2628;
wire _guard2630 = ev00__0state >= 6'd21;
wire _guard2631 = ev00__0state <= 6'd21;
wire _guard2632 = _guard2630 & _guard2631;
wire _guard2633 = ev00__0state >= 6'd21;
wire _guard2634 = ev00__0state <= 6'd21;
wire _guard2635 = _guard2633 & _guard2634;
wire _guard2636 = ev00__0_0;
wire _guard2637 = ev00__0state >= 6'd1;
wire _guard2638 = ev00__0state <= 6'd0;
wire _guard2639 = _guard2637 & _guard2638;
wire _guard2640 = _guard2636 | _guard2639;
wire _guard2641 = ev00__0_0;
wire _guard2642 = ev00__0state >= 6'd1;
wire _guard2643 = ev00__0state <= 6'd0;
wire _guard2644 = _guard2642 & _guard2643;
wire _guard2645 = _guard2641 | _guard2644;
wire _guard2646 = ev00__0_0;
wire _guard2647 = ev00__0state >= 6'd1;
wire _guard2648 = ev00__0state <= 6'd0;
wire _guard2649 = _guard2647 & _guard2648;
wire _guard2650 = _guard2646 | _guard2649;
wire _guard2651 = ev00__0_0;
wire _guard2652 = ev00__0state >= 6'd1;
wire _guard2653 = ev00__0state <= 6'd0;
wire _guard2654 = _guard2652 & _guard2653;
wire _guard2655 = _guard2651 | _guard2654;
wire _guard2656 = ev00__0state >= 6'd44;
wire _guard2657 = ev00__0state <= 6'd44;
wire _guard2658 = _guard2656 & _guard2657;
wire _guard2659 = ev00__0state >= 6'd6;
wire _guard2660 = ev00__0state <= 6'd6;
wire _guard2661 = _guard2659 & _guard2660;
wire _guard2662 = ev00__0_0;
wire _guard2663 = ev00__0state >= 6'd1;
wire _guard2664 = ev00__0state <= 6'd51;
wire _guard2665 = _guard2663 & _guard2664;
wire _guard2666 = _guard2662 | _guard2665;
wire _guard2667 = ev00__0_0;
wire _guard2668 = ev00__0state >= 6'd1;
wire _guard2669 = ev00__0state <= 6'd51;
wire _guard2670 = _guard2668 & _guard2669;
wire _guard2671 = _guard2667 | _guard2670;
wire _guard2672 = ev00__0_0;
wire _guard2673 = ev00__0state >= 6'd1;
wire _guard2674 = ev00__0state <= 6'd51;
wire _guard2675 = _guard2673 & _guard2674;
wire _guard2676 = _guard2672 | _guard2675;
wire _guard2677 = ev00__0_0;
wire _guard2678 = ev00__0state >= 6'd1;
wire _guard2679 = ev00__0state <= 6'd51;
wire _guard2680 = _guard2678 & _guard2679;
wire _guard2681 = _guard2677 | _guard2680;
wire _guard2682 = ev00__0_0;
wire _guard2683 = ev00__0state >= 6'd1;
wire _guard2684 = ev00__0state <= 6'd51;
wire _guard2685 = _guard2683 & _guard2684;
wire _guard2686 = _guard2682 | _guard2685;
wire _guard2687 = ev00__0_0;
wire _guard2688 = ev00__0state >= 6'd1;
wire _guard2689 = ev00__0state <= 6'd51;
wire _guard2690 = _guard2688 & _guard2689;
wire _guard2691 = _guard2687 | _guard2690;
wire _guard2692 = ev00__0_0;
wire _guard2693 = ev00__0state >= 6'd1;
wire _guard2694 = ev00__0state <= 6'd51;
wire _guard2695 = _guard2693 & _guard2694;
wire _guard2696 = _guard2692 | _guard2695;
wire _guard2697 = ev00__0_0;
wire _guard2698 = ev00__0state >= 6'd1;
wire _guard2699 = ev00__0state <= 6'd51;
wire _guard2700 = _guard2698 & _guard2699;
wire _guard2701 = _guard2697 | _guard2700;
wire _guard2702 = ev00__0_0;
wire _guard2703 = ev00__0state >= 6'd1;
wire _guard2704 = ev00__0state <= 6'd51;
wire _guard2705 = _guard2703 & _guard2704;
wire _guard2706 = _guard2702 | _guard2705;
wire _guard2707 = ev00__0_0;
wire _guard2708 = ev00__0state >= 6'd1;
wire _guard2709 = ev00__0state <= 6'd51;
wire _guard2710 = _guard2708 & _guard2709;
wire _guard2711 = _guard2707 | _guard2710;
wire _guard2712 = ev00__0_0;
wire _guard2713 = ev00__0state >= 6'd1;
wire _guard2714 = ev00__0state <= 6'd51;
wire _guard2715 = _guard2713 & _guard2714;
wire _guard2716 = _guard2712 | _guard2715;
wire _guard2717 = ev00__0_0;
wire _guard2718 = ev00__0state >= 6'd1;
wire _guard2719 = ev00__0state <= 6'd51;
wire _guard2720 = _guard2718 & _guard2719;
wire _guard2721 = _guard2717 | _guard2720;
wire _guard2722 = ev00__0_0;
wire _guard2723 = ev00__0state >= 6'd1;
wire _guard2724 = ev00__0state <= 6'd51;
wire _guard2725 = _guard2723 & _guard2724;
wire _guard2726 = _guard2722 | _guard2725;
wire _guard2727 = ev00__0_0;
wire _guard2728 = ev00__0state >= 6'd1;
wire _guard2729 = ev00__0state <= 6'd51;
wire _guard2730 = _guard2728 & _guard2729;
wire _guard2731 = _guard2727 | _guard2730;
wire _guard2732 = ev00__0_0;
wire _guard2733 = ev00__0state >= 6'd1;
wire _guard2734 = ev00__0state <= 6'd51;
wire _guard2735 = _guard2733 & _guard2734;
wire _guard2736 = _guard2732 | _guard2735;
wire _guard2737 = ev00__0_0;
wire _guard2738 = ev00__0state >= 6'd1;
wire _guard2739 = ev00__0state <= 6'd51;
wire _guard2740 = _guard2738 & _guard2739;
wire _guard2741 = _guard2737 | _guard2740;
wire _guard2742 = ev00__0state >= 6'd30;
wire _guard2743 = ev00__0state <= 6'd30;
wire _guard2744 = _guard2742 & _guard2743;
wire _guard2745 = ev00__0state >= 6'd30;
wire _guard2746 = ev00__0state <= 6'd30;
wire _guard2747 = _guard2745 & _guard2746;
wire _guard2748 = ev00__0state >= 6'd30;
wire _guard2749 = ev00__0state <= 6'd30;
wire _guard2750 = _guard2748 & _guard2749;
wire _guard2751 = ev00__0state >= 6'd30;
wire _guard2752 = ev00__0state <= 6'd30;
wire _guard2753 = _guard2751 & _guard2752;
wire _guard2754 = ev00__0state >= 6'd18;
wire _guard2755 = ev00__0state <= 6'd18;
wire _guard2756 = _guard2754 & _guard2755;
wire _guard2757 = ev00__0state >= 6'd18;
wire _guard2758 = ev00__0state <= 6'd18;
wire _guard2759 = _guard2757 & _guard2758;
wire _guard2760 = ev00__0state >= 6'd18;
wire _guard2761 = ev00__0state <= 6'd18;
wire _guard2762 = _guard2760 & _guard2761;
wire _guard2763 = ev00__0state >= 6'd18;
wire _guard2764 = ev00__0state <= 6'd18;
wire _guard2765 = _guard2763 & _guard2764;
wire _guard2766 = ev00__0_0;
wire _guard2767 = ev00__0state >= 6'd1;
wire _guard2768 = ev00__0state <= 6'd0;
wire _guard2769 = _guard2767 & _guard2768;
wire _guard2770 = _guard2766 | _guard2769;
wire _guard2771 = ev00__0state >= 6'd8;
wire _guard2772 = ev00__0state <= 6'd8;
wire _guard2773 = _guard2771 & _guard2772;
wire _guard2774 = _guard2770 | _guard2773;
wire _guard2775 = ev00__0state >= 6'd13;
wire _guard2776 = ev00__0state <= 6'd13;
wire _guard2777 = _guard2775 & _guard2776;
wire _guard2778 = _guard2774 | _guard2777;
wire _guard2779 = ev00__0state >= 6'd21;
wire _guard2780 = ev00__0state <= 6'd21;
wire _guard2781 = _guard2779 & _guard2780;
wire _guard2782 = _guard2778 | _guard2781;
wire _guard2783 = ev00__0state >= 6'd26;
wire _guard2784 = ev00__0state <= 6'd26;
wire _guard2785 = _guard2783 & _guard2784;
wire _guard2786 = _guard2782 | _guard2785;
wire _guard2787 = ev00__0state >= 6'd34;
wire _guard2788 = ev00__0state <= 6'd34;
wire _guard2789 = _guard2787 & _guard2788;
wire _guard2790 = _guard2786 | _guard2789;
wire _guard2791 = ev00__0state >= 6'd39;
wire _guard2792 = ev00__0state <= 6'd39;
wire _guard2793 = _guard2791 & _guard2792;
wire _guard2794 = _guard2790 | _guard2793;
wire _guard2795 = ev00__0state >= 6'd47;
wire _guard2796 = ev00__0state <= 6'd47;
wire _guard2797 = _guard2795 & _guard2796;
wire _guard2798 = _guard2794 | _guard2797;
wire _guard2799 = ev00__0state >= 6'd26;
wire _guard2800 = ev00__0state <= 6'd26;
wire _guard2801 = _guard2799 & _guard2800;
wire _guard2802 = ev00__0state >= 6'd8;
wire _guard2803 = ev00__0state <= 6'd8;
wire _guard2804 = _guard2802 & _guard2803;
wire _guard2805 = ev00__0state >= 6'd13;
wire _guard2806 = ev00__0state <= 6'd13;
wire _guard2807 = _guard2805 & _guard2806;
wire _guard2808 = ev00__0state >= 6'd34;
wire _guard2809 = ev00__0state <= 6'd34;
wire _guard2810 = _guard2808 & _guard2809;
wire _guard2811 = ev00__0state >= 6'd21;
wire _guard2812 = ev00__0state <= 6'd21;
wire _guard2813 = _guard2811 & _guard2812;
wire _guard2814 = ev00__0_0;
wire _guard2815 = ev00__0state >= 6'd1;
wire _guard2816 = ev00__0state <= 6'd0;
wire _guard2817 = _guard2815 & _guard2816;
wire _guard2818 = _guard2814 | _guard2817;
wire _guard2819 = ev00__0state >= 6'd39;
wire _guard2820 = ev00__0state <= 6'd39;
wire _guard2821 = _guard2819 & _guard2820;
wire _guard2822 = ev00__0state >= 6'd47;
wire _guard2823 = ev00__0state <= 6'd47;
wire _guard2824 = _guard2822 & _guard2823;
wire _guard2825 = ev00__0_0;
wire _guard2826 = ev00__0state >= 6'd1;
wire _guard2827 = ev00__0state <= 6'd0;
wire _guard2828 = _guard2826 & _guard2827;
wire _guard2829 = _guard2825 | _guard2828;
wire _guard2830 = ev00__0_0;
wire _guard2831 = ev00__0state >= 6'd1;
wire _guard2832 = ev00__0state <= 6'd0;
wire _guard2833 = _guard2831 & _guard2832;
wire _guard2834 = _guard2830 | _guard2833;
wire _guard2835 = ev00__0_0;
wire _guard2836 = ev00__0state >= 6'd1;
wire _guard2837 = ev00__0state <= 6'd0;
wire _guard2838 = _guard2836 & _guard2837;
wire _guard2839 = _guard2835 | _guard2838;
wire _guard2840 = ev00__0_0;
wire _guard2841 = ev00__0state >= 6'd1;
wire _guard2842 = ev00__0state <= 6'd0;
wire _guard2843 = _guard2841 & _guard2842;
wire _guard2844 = _guard2840 | _guard2843;
wire _guard2845 = ev00__0state >= 6'd51;
wire _guard2846 = ev00__0state <= 6'd51;
wire _guard2847 = _guard2845 & _guard2846;
wire _guard2848 = ev00__0state >= 6'd12;
wire _guard2849 = ev00__0state <= 6'd12;
wire _guard2850 = _guard2848 & _guard2849;
wire _guard2851 = ev00__0state >= 6'd26;
wire _guard2852 = ev00__0state <= 6'd26;
wire _guard2853 = _guard2851 & _guard2852;
wire _guard2854 = ev00__0state >= 6'd26;
wire _guard2855 = ev00__0state <= 6'd26;
wire _guard2856 = _guard2854 & _guard2855;
wire _guard2857 = ev00__0state >= 6'd26;
wire _guard2858 = ev00__0state <= 6'd26;
wire _guard2859 = _guard2857 & _guard2858;
wire _guard2860 = ev00__0state >= 6'd26;
wire _guard2861 = ev00__0state <= 6'd26;
wire _guard2862 = _guard2860 & _guard2861;
wire _guard2863 = ev00__0state >= 6'd38;
wire _guard2864 = ev00__0state <= 6'd38;
wire _guard2865 = _guard2863 & _guard2864;
wire _guard2866 = ev00__0state >= 6'd38;
wire _guard2867 = ev00__0state <= 6'd38;
wire _guard2868 = _guard2866 & _guard2867;
wire _guard2869 = ev00__0state >= 6'd38;
wire _guard2870 = ev00__0state <= 6'd38;
wire _guard2871 = _guard2869 & _guard2870;
wire _guard2872 = ev00__0state >= 6'd38;
wire _guard2873 = ev00__0state <= 6'd38;
wire _guard2874 = _guard2872 & _guard2873;
wire _guard2875 = ev00__0state >= 6'd38;
wire _guard2876 = ev00__0state <= 6'd38;
wire _guard2877 = _guard2875 & _guard2876;
wire _guard2878 = ev00__0state >= 6'd38;
wire _guard2879 = ev00__0state <= 6'd38;
wire _guard2880 = _guard2878 & _guard2879;
wire _guard2881 = ev00__0state >= 6'd38;
wire _guard2882 = ev00__0state <= 6'd38;
wire _guard2883 = _guard2881 & _guard2882;
wire _guard2884 = ev00__0state >= 6'd38;
wire _guard2885 = ev00__0state <= 6'd38;
wire _guard2886 = _guard2884 & _guard2885;
wire _guard2887 = ev00__0state >= 6'd38;
wire _guard2888 = ev00__0state <= 6'd38;
wire _guard2889 = _guard2887 & _guard2888;
wire _guard2890 = ev00__0state >= 6'd38;
wire _guard2891 = ev00__0state <= 6'd38;
wire _guard2892 = _guard2890 & _guard2891;
wire _guard2893 = ev00__0state >= 6'd38;
wire _guard2894 = ev00__0state <= 6'd38;
wire _guard2895 = _guard2893 & _guard2894;
wire _guard2896 = ev00__0state >= 6'd38;
wire _guard2897 = ev00__0state <= 6'd38;
wire _guard2898 = _guard2896 & _guard2897;
wire _guard2899 = ev00__0state >= 6'd38;
wire _guard2900 = ev00__0state <= 6'd38;
wire _guard2901 = _guard2899 & _guard2900;
wire _guard2902 = ev00__0state >= 6'd38;
wire _guard2903 = ev00__0state <= 6'd38;
wire _guard2904 = _guard2902 & _guard2903;
wire _guard2905 = ev00__0state >= 6'd38;
wire _guard2906 = ev00__0state <= 6'd38;
wire _guard2907 = _guard2905 & _guard2906;
wire _guard2908 = ev00__0state >= 6'd38;
wire _guard2909 = ev00__0state <= 6'd38;
wire _guard2910 = _guard2908 & _guard2909;
wire _guard2911 = ev00__0state >= 6'd38;
wire _guard2912 = ev00__0state <= 6'd38;
wire _guard2913 = _guard2911 & _guard2912;
wire _guard2914 = ev00__0state >= 6'd38;
wire _guard2915 = ev00__0state <= 6'd38;
wire _guard2916 = _guard2914 & _guard2915;
wire _guard2917 = ev00__0state >= 6'd38;
wire _guard2918 = ev00__0state <= 6'd38;
wire _guard2919 = _guard2917 & _guard2918;
wire _guard2920 = ev00__0state >= 6'd38;
wire _guard2921 = ev00__0state <= 6'd38;
wire _guard2922 = _guard2920 & _guard2921;
wire _guard2923 = ev00__0state >= 6'd38;
wire _guard2924 = ev00__0state <= 6'd38;
wire _guard2925 = _guard2923 & _guard2924;
wire _guard2926 = ev00__0state >= 6'd38;
wire _guard2927 = ev00__0state <= 6'd38;
wire _guard2928 = _guard2926 & _guard2927;
wire _guard2929 = ev00__0state >= 6'd38;
wire _guard2930 = ev00__0state <= 6'd38;
wire _guard2931 = _guard2929 & _guard2930;
wire _guard2932 = ev00__0state >= 6'd38;
wire _guard2933 = ev00__0state <= 6'd38;
wire _guard2934 = _guard2932 & _guard2933;
wire _guard2935 = ev00__0state >= 6'd38;
wire _guard2936 = ev00__0state <= 6'd38;
wire _guard2937 = _guard2935 & _guard2936;
wire _guard2938 = ev00__0state >= 6'd38;
wire _guard2939 = ev00__0state <= 6'd38;
wire _guard2940 = _guard2938 & _guard2939;
wire _guard2941 = ev00__0state >= 6'd38;
wire _guard2942 = ev00__0state <= 6'd38;
wire _guard2943 = _guard2941 & _guard2942;
wire _guard2944 = ev00__0state >= 6'd38;
wire _guard2945 = ev00__0state <= 6'd38;
wire _guard2946 = _guard2944 & _guard2945;
wire _guard2947 = ev00__0state >= 6'd38;
wire _guard2948 = ev00__0state <= 6'd38;
wire _guard2949 = _guard2947 & _guard2948;
wire _guard2950 = ev00__0state >= 6'd38;
wire _guard2951 = ev00__0state <= 6'd38;
wire _guard2952 = _guard2950 & _guard2951;
wire _guard2953 = ev00__0state >= 6'd38;
wire _guard2954 = ev00__0state <= 6'd38;
wire _guard2955 = _guard2953 & _guard2954;
wire _guard2956 = ev00__0state >= 6'd38;
wire _guard2957 = ev00__0state <= 6'd38;
wire _guard2958 = _guard2956 & _guard2957;
wire _guard2959 = ev00__0state >= 6'd38;
wire _guard2960 = ev00__0state <= 6'd38;
wire _guard2961 = _guard2959 & _guard2960;
wire _guard2962 = ev00__0state >= 6'd13;
wire _guard2963 = ev00__0state <= 6'd13;
wire _guard2964 = _guard2962 & _guard2963;
wire _guard2965 = ev00__0state >= 6'd26;
wire _guard2966 = ev00__0state <= 6'd26;
wire _guard2967 = _guard2965 & _guard2966;
wire _guard2968 = ev00__0state >= 6'd39;
wire _guard2969 = ev00__0state <= 6'd39;
wire _guard2970 = _guard2968 & _guard2969;
wire _guard2971 = ev00__0_0;
wire _guard2972 = ev00__0state >= 6'd1;
wire _guard2973 = ev00__0state <= 6'd0;
wire _guard2974 = _guard2972 & _guard2973;
wire _guard2975 = _guard2971 | _guard2974;
wire _guard2976 = ev00__0state >= 6'd5;
wire _guard2977 = ev00__0state <= 6'd5;
wire _guard2978 = _guard2976 & _guard2977;
wire _guard2979 = _guard2975 | _guard2978;
wire _guard2980 = ev00__0state >= 6'd13;
wire _guard2981 = ev00__0state <= 6'd13;
wire _guard2982 = _guard2980 & _guard2981;
wire _guard2983 = _guard2979 | _guard2982;
wire _guard2984 = ev00__0state >= 6'd18;
wire _guard2985 = ev00__0state <= 6'd18;
wire _guard2986 = _guard2984 & _guard2985;
wire _guard2987 = _guard2983 | _guard2986;
wire _guard2988 = ev00__0state >= 6'd26;
wire _guard2989 = ev00__0state <= 6'd26;
wire _guard2990 = _guard2988 & _guard2989;
wire _guard2991 = _guard2987 | _guard2990;
wire _guard2992 = ev00__0state >= 6'd31;
wire _guard2993 = ev00__0state <= 6'd31;
wire _guard2994 = _guard2992 & _guard2993;
wire _guard2995 = _guard2991 | _guard2994;
wire _guard2996 = ev00__0state >= 6'd39;
wire _guard2997 = ev00__0state <= 6'd39;
wire _guard2998 = _guard2996 & _guard2997;
wire _guard2999 = _guard2995 | _guard2998;
wire _guard3000 = ev00__0state >= 6'd44;
wire _guard3001 = ev00__0state <= 6'd44;
wire _guard3002 = _guard3000 & _guard3001;
wire _guard3003 = _guard2999 | _guard3002;
wire _guard3004 = ev00__0state >= 6'd44;
wire _guard3005 = ev00__0state <= 6'd44;
wire _guard3006 = _guard3004 & _guard3005;
wire _guard3007 = ev00__0state >= 6'd13;
wire _guard3008 = ev00__0state <= 6'd13;
wire _guard3009 = _guard3007 & _guard3008;
wire _guard3010 = ev00__0state >= 6'd5;
wire _guard3011 = ev00__0state <= 6'd5;
wire _guard3012 = _guard3010 & _guard3011;
wire _guard3013 = ev00__0_0;
wire _guard3014 = ev00__0state >= 6'd1;
wire _guard3015 = ev00__0state <= 6'd0;
wire _guard3016 = _guard3014 & _guard3015;
wire _guard3017 = _guard3013 | _guard3016;
wire _guard3018 = ev00__0state >= 6'd39;
wire _guard3019 = ev00__0state <= 6'd39;
wire _guard3020 = _guard3018 & _guard3019;
wire _guard3021 = ev00__0state >= 6'd18;
wire _guard3022 = ev00__0state <= 6'd18;
wire _guard3023 = _guard3021 & _guard3022;
wire _guard3024 = ev00__0state >= 6'd31;
wire _guard3025 = ev00__0state <= 6'd31;
wire _guard3026 = _guard3024 & _guard3025;
wire _guard3027 = ev00__0state >= 6'd26;
wire _guard3028 = ev00__0state <= 6'd26;
wire _guard3029 = _guard3027 & _guard3028;
wire _guard3030 = ev00__0state >= 6'd31;
wire _guard3031 = ev00__0state <= 6'd31;
wire _guard3032 = _guard3030 & _guard3031;
wire _guard3033 = ev00__0state >= 6'd31;
wire _guard3034 = ev00__0state <= 6'd31;
wire _guard3035 = _guard3033 & _guard3034;
wire _guard3036 = ev00__0state >= 6'd31;
wire _guard3037 = ev00__0state <= 6'd31;
wire _guard3038 = _guard3036 & _guard3037;
wire _guard3039 = ev00__0state >= 6'd31;
wire _guard3040 = ev00__0state <= 6'd31;
wire _guard3041 = _guard3039 & _guard3040;
wire _guard3042 = ev00__0state >= 6'd7;
wire _guard3043 = ev00__0state <= 6'd7;
wire _guard3044 = _guard3042 & _guard3043;
wire _guard3045 = ev00__0state >= 6'd7;
wire _guard3046 = ev00__0state <= 6'd7;
wire _guard3047 = _guard3045 & _guard3046;
wire _guard3048 = ev00__0state >= 6'd7;
wire _guard3049 = ev00__0state <= 6'd7;
wire _guard3050 = _guard3048 & _guard3049;
wire _guard3051 = ev00__0state >= 6'd7;
wire _guard3052 = ev00__0state <= 6'd7;
wire _guard3053 = _guard3051 & _guard3052;
wire _guard3054 = ev00__0state >= 6'd20;
wire _guard3055 = ev00__0state <= 6'd20;
wire _guard3056 = _guard3054 & _guard3055;
wire _guard3057 = ev00__0state >= 6'd20;
wire _guard3058 = ev00__0state <= 6'd20;
wire _guard3059 = _guard3057 & _guard3058;
wire _guard3060 = ev00__0state >= 6'd20;
wire _guard3061 = ev00__0state <= 6'd20;
wire _guard3062 = _guard3060 & _guard3061;
wire _guard3063 = ev00__0state >= 6'd20;
wire _guard3064 = ev00__0state <= 6'd20;
wire _guard3065 = _guard3063 & _guard3064;
wire _guard3066 = ev00__0state >= 6'd30;
wire _guard3067 = ev00__0state <= 6'd30;
wire _guard3068 = _guard3066 & _guard3067;
wire _guard3069 = ev00__0state >= 6'd38;
wire _guard3070 = ev00__0state <= 6'd38;
wire _guard3071 = _guard3069 & _guard3070;
wire _guard3072 = ev00__0state >= 6'd35;
wire _guard3073 = ev00__0state <= 6'd35;
wire _guard3074 = _guard3072 & _guard3073;
wire _guard3075 = ev00__0state >= 6'd35;
wire _guard3076 = ev00__0state <= 6'd35;
wire _guard3077 = _guard3075 & _guard3076;
wire _guard3078 = ev00__0state >= 6'd35;
wire _guard3079 = ev00__0state <= 6'd35;
wire _guard3080 = _guard3078 & _guard3079;
wire _guard3081 = ev00__0state >= 6'd35;
wire _guard3082 = ev00__0state <= 6'd35;
wire _guard3083 = _guard3081 & _guard3082;
wire _guard3084 = ev00__0_0;
wire _guard3085 = ev00__0state >= 6'd1;
wire _guard3086 = ev00__0state <= 6'd0;
wire _guard3087 = _guard3085 & _guard3086;
wire _guard3088 = _guard3084 | _guard3087;
wire _guard3089 = ev00__0_0;
wire _guard3090 = ev00__0state >= 6'd1;
wire _guard3091 = ev00__0state <= 6'd0;
wire _guard3092 = _guard3090 & _guard3091;
wire _guard3093 = _guard3089 | _guard3092;
wire _guard3094 = ev00__0_0;
wire _guard3095 = ev00__0state >= 6'd1;
wire _guard3096 = ev00__0state <= 6'd0;
wire _guard3097 = _guard3095 & _guard3096;
wire _guard3098 = _guard3094 | _guard3097;
wire _guard3099 = ev00__0_0;
wire _guard3100 = ev00__0state >= 6'd1;
wire _guard3101 = ev00__0state <= 6'd0;
wire _guard3102 = _guard3100 & _guard3101;
wire _guard3103 = _guard3099 | _guard3102;
wire _guard3104 = ev00__0state >= 6'd25;
wire _guard3105 = ev00__0state <= 6'd25;
wire _guard3106 = _guard3104 & _guard3105;
wire _guard3107 = ev00__0state >= 6'd36;
wire _guard3108 = ev00__0state <= 6'd36;
wire _guard3109 = _guard3107 & _guard3108;
wire _guard3110 = ev00__0state >= 6'd36;
wire _guard3111 = ev00__0state <= 6'd36;
wire _guard3112 = _guard3110 & _guard3111;
wire _guard3113 = ev00__0state >= 6'd36;
wire _guard3114 = ev00__0state <= 6'd36;
wire _guard3115 = _guard3113 & _guard3114;
wire _guard3116 = ev00__0state >= 6'd36;
wire _guard3117 = ev00__0state <= 6'd36;
wire _guard3118 = _guard3116 & _guard3117;
wire _guard3119 = ev00__0state >= 6'd51;
wire _guard3120 = ev00__0state <= 6'd51;
wire _guard3121 = _guard3119 & _guard3120;
wire _guard3122 = ev00__0state >= 6'd25;
wire _guard3123 = ev00__0state <= 6'd25;
wire _guard3124 = _guard3122 & _guard3123;
wire _guard3125 = ev00__0state >= 6'd51;
wire _guard3126 = ev00__0state <= 6'd51;
wire _guard3127 = _guard3125 & _guard3126;
wire _guard3128 = ev00__0state >= 6'd38;
wire _guard3129 = ev00__0state <= 6'd38;
wire _guard3130 = _guard3128 & _guard3129;
wire _guard3131 = ev00__0state >= 6'd12;
wire _guard3132 = ev00__0state <= 6'd12;
wire _guard3133 = _guard3131 & _guard3132;
wire _guard3134 = ev00__0state >= 6'd12;
wire _guard3135 = ev00__0state <= 6'd12;
wire _guard3136 = _guard3134 & _guard3135;
wire _guard3137 = ev00__0state >= 6'd38;
wire _guard3138 = ev00__0state <= 6'd38;
wire _guard3139 = _guard3137 & _guard3138;
wire _guard3140 = ev00__0state >= 6'd25;
wire _guard3141 = ev00__0state <= 6'd25;
wire _guard3142 = _guard3140 & _guard3141;
wire _guard3143 = ev00__0state >= 6'd51;
wire _guard3144 = ev00__0state <= 6'd51;
wire _guard3145 = _guard3143 & _guard3144;
wire _guard3146 = ev00__0state >= 6'd12;
wire _guard3147 = ev00__0state <= 6'd12;
wire _guard3148 = _guard3146 & _guard3147;
wire _guard3149 = ev00__0state >= 6'd38;
wire _guard3150 = ev00__0state <= 6'd38;
wire _guard3151 = _guard3149 & _guard3150;
wire _guard3152 = ev00__0state >= 6'd25;
wire _guard3153 = ev00__0state <= 6'd25;
wire _guard3154 = _guard3152 & _guard3153;
wire _guard3155 = ev00__0state >= 6'd51;
wire _guard3156 = ev00__0state <= 6'd51;
wire _guard3157 = _guard3155 & _guard3156;
wire _guard3158 = ev00__0state >= 6'd38;
wire _guard3159 = ev00__0state <= 6'd38;
wire _guard3160 = _guard3158 & _guard3159;
wire _guard3161 = ev00__0state >= 6'd25;
wire _guard3162 = ev00__0state <= 6'd25;
wire _guard3163 = _guard3161 & _guard3162;
wire _guard3164 = ev00__0state >= 6'd51;
wire _guard3165 = ev00__0state <= 6'd51;
wire _guard3166 = _guard3164 & _guard3165;
wire _guard3167 = ev00__0state >= 6'd12;
wire _guard3168 = ev00__0state <= 6'd12;
wire _guard3169 = _guard3167 & _guard3168;
wire _guard3170 = ev00__0state >= 6'd38;
wire _guard3171 = ev00__0state <= 6'd38;
wire _guard3172 = _guard3170 & _guard3171;
wire _guard3173 = ev00__0state >= 6'd25;
wire _guard3174 = ev00__0state <= 6'd25;
wire _guard3175 = _guard3173 & _guard3174;
wire _guard3176 = ev00__0state >= 6'd51;
wire _guard3177 = ev00__0state <= 6'd51;
wire _guard3178 = _guard3176 & _guard3177;
wire _guard3179 = ev00__0state >= 6'd12;
wire _guard3180 = ev00__0state <= 6'd12;
wire _guard3181 = _guard3179 & _guard3180;
wire _guard3182 = ev00__0state >= 6'd38;
wire _guard3183 = ev00__0state <= 6'd38;
wire _guard3184 = _guard3182 & _guard3183;
wire _guard3185 = ev00__0state >= 6'd51;
wire _guard3186 = ev00__0state <= 6'd51;
wire _guard3187 = _guard3185 & _guard3186;
wire _guard3188 = ev00__0state >= 6'd25;
wire _guard3189 = ev00__0state <= 6'd25;
wire _guard3190 = _guard3188 & _guard3189;
wire _guard3191 = ev00__0state >= 6'd12;
wire _guard3192 = ev00__0state <= 6'd12;
wire _guard3193 = _guard3191 & _guard3192;
wire _guard3194 = ev00__0state >= 6'd38;
wire _guard3195 = ev00__0state <= 6'd38;
wire _guard3196 = _guard3194 & _guard3195;
wire _guard3197 = ev00__0state >= 6'd25;
wire _guard3198 = ev00__0state <= 6'd25;
wire _guard3199 = _guard3197 & _guard3198;
wire _guard3200 = ev00__0state >= 6'd51;
wire _guard3201 = ev00__0state <= 6'd51;
wire _guard3202 = _guard3200 & _guard3201;
wire _guard3203 = ev00__0state >= 6'd12;
wire _guard3204 = ev00__0state <= 6'd12;
wire _guard3205 = _guard3203 & _guard3204;
wire _guard3206 = ev00__0state >= 6'd38;
wire _guard3207 = ev00__0state <= 6'd38;
wire _guard3208 = _guard3206 & _guard3207;
wire _guard3209 = ev00__0state >= 6'd25;
wire _guard3210 = ev00__0state <= 6'd25;
wire _guard3211 = _guard3209 & _guard3210;
wire _guard3212 = ev00__0state >= 6'd51;
wire _guard3213 = ev00__0state <= 6'd51;
wire _guard3214 = _guard3212 & _guard3213;
wire _guard3215 = ev00__0state >= 6'd12;
wire _guard3216 = ev00__0state <= 6'd12;
wire _guard3217 = _guard3215 & _guard3216;
wire _guard3218 = ev00__0state >= 6'd38;
wire _guard3219 = ev00__0state <= 6'd38;
wire _guard3220 = _guard3218 & _guard3219;
wire _guard3221 = ev00__0state >= 6'd25;
wire _guard3222 = ev00__0state <= 6'd25;
wire _guard3223 = _guard3221 & _guard3222;
wire _guard3224 = ev00__0state >= 6'd51;
wire _guard3225 = ev00__0state <= 6'd51;
wire _guard3226 = _guard3224 & _guard3225;
wire _guard3227 = ev00__0state >= 6'd12;
wire _guard3228 = ev00__0state <= 6'd12;
wire _guard3229 = _guard3227 & _guard3228;
wire _guard3230 = ev00__0state >= 6'd38;
wire _guard3231 = ev00__0state <= 6'd38;
wire _guard3232 = _guard3230 & _guard3231;
wire _guard3233 = ev00__0state >= 6'd25;
wire _guard3234 = ev00__0state <= 6'd25;
wire _guard3235 = _guard3233 & _guard3234;
wire _guard3236 = ev00__0state >= 6'd51;
wire _guard3237 = ev00__0state <= 6'd51;
wire _guard3238 = _guard3236 & _guard3237;
wire _guard3239 = ev00__0state >= 6'd12;
wire _guard3240 = ev00__0state <= 6'd12;
wire _guard3241 = _guard3239 & _guard3240;
wire _guard3242 = ev00__0state >= 6'd25;
wire _guard3243 = ev00__0state <= 6'd25;
wire _guard3244 = _guard3242 & _guard3243;
wire _guard3245 = ev00__0state >= 6'd51;
wire _guard3246 = ev00__0state <= 6'd51;
wire _guard3247 = _guard3245 & _guard3246;
wire _guard3248 = ev00__0state >= 6'd38;
wire _guard3249 = ev00__0state <= 6'd38;
wire _guard3250 = _guard3248 & _guard3249;
wire _guard3251 = ev00__0state >= 6'd12;
wire _guard3252 = ev00__0state <= 6'd12;
wire _guard3253 = _guard3251 & _guard3252;
wire _guard3254 = ev00__0state >= 6'd25;
wire _guard3255 = ev00__0state <= 6'd25;
wire _guard3256 = _guard3254 & _guard3255;
wire _guard3257 = ev00__0state >= 6'd51;
wire _guard3258 = ev00__0state <= 6'd51;
wire _guard3259 = _guard3257 & _guard3258;
wire _guard3260 = ev00__0state >= 6'd38;
wire _guard3261 = ev00__0state <= 6'd38;
wire _guard3262 = _guard3260 & _guard3261;
wire _guard3263 = ev00__0state >= 6'd12;
wire _guard3264 = ev00__0state <= 6'd12;
wire _guard3265 = _guard3263 & _guard3264;
wire _guard3266 = ev00__0state >= 6'd38;
wire _guard3267 = ev00__0state <= 6'd38;
wire _guard3268 = _guard3266 & _guard3267;
wire _guard3269 = ev00__0state >= 6'd12;
wire _guard3270 = ev00__0state <= 6'd12;
wire _guard3271 = _guard3269 & _guard3270;
wire _guard3272 = ev00__0state >= 6'd25;
wire _guard3273 = ev00__0state <= 6'd25;
wire _guard3274 = _guard3272 & _guard3273;
wire _guard3275 = ev00__0state >= 6'd51;
wire _guard3276 = ev00__0state <= 6'd51;
wire _guard3277 = _guard3275 & _guard3276;
wire _guard3278 = ev00__0state >= 6'd38;
wire _guard3279 = ev00__0state <= 6'd38;
wire _guard3280 = _guard3278 & _guard3279;
wire _guard3281 = ev00__0state >= 6'd25;
wire _guard3282 = ev00__0state <= 6'd25;
wire _guard3283 = _guard3281 & _guard3282;
wire _guard3284 = ev00__0state >= 6'd51;
wire _guard3285 = ev00__0state <= 6'd51;
wire _guard3286 = _guard3284 & _guard3285;
wire _guard3287 = ev00__0state >= 6'd12;
wire _guard3288 = ev00__0state <= 6'd12;
wire _guard3289 = _guard3287 & _guard3288;
wire _guard3290 = ev00__0state >= 6'd38;
wire _guard3291 = ev00__0state <= 6'd38;
wire _guard3292 = _guard3290 & _guard3291;
wire _guard3293 = ev00__0state >= 6'd12;
wire _guard3294 = ev00__0state <= 6'd12;
wire _guard3295 = _guard3293 & _guard3294;
wire _guard3296 = ev00__0state >= 6'd25;
wire _guard3297 = ev00__0state <= 6'd25;
wire _guard3298 = _guard3296 & _guard3297;
wire _guard3299 = ev00__0state >= 6'd51;
wire _guard3300 = ev00__0state <= 6'd51;
wire _guard3301 = _guard3299 & _guard3300;
wire _guard3302 = ev00__0state >= 6'd38;
wire _guard3303 = ev00__0state <= 6'd38;
wire _guard3304 = _guard3302 & _guard3303;
wire _guard3305 = ev00__0state >= 6'd51;
wire _guard3306 = ev00__0state <= 6'd51;
wire _guard3307 = _guard3305 & _guard3306;
wire _guard3308 = ev00__0state >= 6'd25;
wire _guard3309 = ev00__0state <= 6'd25;
wire _guard3310 = _guard3308 & _guard3309;
wire _guard3311 = ev00__0state >= 6'd12;
wire _guard3312 = ev00__0state <= 6'd12;
wire _guard3313 = _guard3311 & _guard3312;
wire _guard3314 = ev00__0state >= 6'd38;
wire _guard3315 = ev00__0state <= 6'd38;
wire _guard3316 = _guard3314 & _guard3315;
wire _guard3317 = ev00__0state >= 6'd25;
wire _guard3318 = ev00__0state <= 6'd25;
wire _guard3319 = _guard3317 & _guard3318;
wire _guard3320 = ev00__0state >= 6'd51;
wire _guard3321 = ev00__0state <= 6'd51;
wire _guard3322 = _guard3320 & _guard3321;
wire _guard3323 = ev00__0state >= 6'd12;
wire _guard3324 = ev00__0state <= 6'd12;
wire _guard3325 = _guard3323 & _guard3324;
wire _guard3326 = ev00__0state >= 6'd38;
wire _guard3327 = ev00__0state <= 6'd38;
wire _guard3328 = _guard3326 & _guard3327;
wire _guard3329 = ev00__0state >= 6'd25;
wire _guard3330 = ev00__0state <= 6'd25;
wire _guard3331 = _guard3329 & _guard3330;
wire _guard3332 = ev00__0state >= 6'd51;
wire _guard3333 = ev00__0state <= 6'd51;
wire _guard3334 = _guard3332 & _guard3333;
wire _guard3335 = ev00__0state >= 6'd12;
wire _guard3336 = ev00__0state <= 6'd12;
wire _guard3337 = _guard3335 & _guard3336;
wire _guard3338 = ev00__0state >= 6'd38;
wire _guard3339 = ev00__0state <= 6'd38;
wire _guard3340 = _guard3338 & _guard3339;
wire _guard3341 = ev00__0state >= 6'd51;
wire _guard3342 = ev00__0state <= 6'd51;
wire _guard3343 = _guard3341 & _guard3342;
wire _guard3344 = ev00__0state >= 6'd25;
wire _guard3345 = ev00__0state <= 6'd25;
wire _guard3346 = _guard3344 & _guard3345;
wire _guard3347 = ev00__0state >= 6'd12;
wire _guard3348 = ev00__0state <= 6'd12;
wire _guard3349 = _guard3347 & _guard3348;
wire _guard3350 = ev00__0state >= 6'd38;
wire _guard3351 = ev00__0state <= 6'd38;
wire _guard3352 = _guard3350 & _guard3351;
wire _guard3353 = ev00__0state >= 6'd51;
wire _guard3354 = ev00__0state <= 6'd51;
wire _guard3355 = _guard3353 & _guard3354;
wire _guard3356 = ev00__0state >= 6'd25;
wire _guard3357 = ev00__0state <= 6'd25;
wire _guard3358 = _guard3356 & _guard3357;
wire _guard3359 = ev00__0state >= 6'd12;
wire _guard3360 = ev00__0state <= 6'd12;
wire _guard3361 = _guard3359 & _guard3360;
wire _guard3362 = ev00__0state >= 6'd38;
wire _guard3363 = ev00__0state <= 6'd38;
wire _guard3364 = _guard3362 & _guard3363;
wire _guard3365 = ev00__0state >= 6'd25;
wire _guard3366 = ev00__0state <= 6'd25;
wire _guard3367 = _guard3365 & _guard3366;
wire _guard3368 = ev00__0state >= 6'd51;
wire _guard3369 = ev00__0state <= 6'd51;
wire _guard3370 = _guard3368 & _guard3369;
wire _guard3371 = ev00__0state >= 6'd12;
wire _guard3372 = ev00__0state <= 6'd12;
wire _guard3373 = _guard3371 & _guard3372;
wire _guard3374 = ev00__0state >= 6'd38;
wire _guard3375 = ev00__0state <= 6'd38;
wire _guard3376 = _guard3374 & _guard3375;
wire _guard3377 = ev00__0state >= 6'd25;
wire _guard3378 = ev00__0state <= 6'd25;
wire _guard3379 = _guard3377 & _guard3378;
wire _guard3380 = ev00__0state >= 6'd51;
wire _guard3381 = ev00__0state <= 6'd51;
wire _guard3382 = _guard3380 & _guard3381;
wire _guard3383 = ev00__0state >= 6'd12;
wire _guard3384 = ev00__0state <= 6'd12;
wire _guard3385 = _guard3383 & _guard3384;
wire _guard3386 = ev00__0state >= 6'd25;
wire _guard3387 = ev00__0state <= 6'd25;
wire _guard3388 = _guard3386 & _guard3387;
wire _guard3389 = ev00__0state >= 6'd51;
wire _guard3390 = ev00__0state <= 6'd51;
wire _guard3391 = _guard3389 & _guard3390;
wire _guard3392 = ev00__0state >= 6'd38;
wire _guard3393 = ev00__0state <= 6'd38;
wire _guard3394 = _guard3392 & _guard3393;
wire _guard3395 = ev00__0state >= 6'd12;
wire _guard3396 = ev00__0state <= 6'd12;
wire _guard3397 = _guard3395 & _guard3396;
wire _guard3398 = ev00__0state >= 6'd38;
wire _guard3399 = ev00__0state <= 6'd38;
wire _guard3400 = _guard3398 & _guard3399;
wire _guard3401 = ev00__0state >= 6'd25;
wire _guard3402 = ev00__0state <= 6'd25;
wire _guard3403 = _guard3401 & _guard3402;
wire _guard3404 = ev00__0state >= 6'd12;
wire _guard3405 = ev00__0state <= 6'd12;
wire _guard3406 = _guard3404 & _guard3405;
wire _guard3407 = ev00__0state >= 6'd51;
wire _guard3408 = ev00__0state <= 6'd51;
wire _guard3409 = _guard3407 & _guard3408;
wire _guard3410 = ev00__0state >= 6'd38;
wire _guard3411 = ev00__0state <= 6'd38;
wire _guard3412 = _guard3410 & _guard3411;
wire _guard3413 = ev00__0state >= 6'd12;
wire _guard3414 = ev00__0state <= 6'd12;
wire _guard3415 = _guard3413 & _guard3414;
wire _guard3416 = ev00__0state >= 6'd25;
wire _guard3417 = ev00__0state <= 6'd25;
wire _guard3418 = _guard3416 & _guard3417;
wire _guard3419 = ev00__0state >= 6'd51;
wire _guard3420 = ev00__0state <= 6'd51;
wire _guard3421 = _guard3419 & _guard3420;
wire _guard3422 = ev00__0state >= 6'd38;
wire _guard3423 = ev00__0state <= 6'd38;
wire _guard3424 = _guard3422 & _guard3423;
wire _guard3425 = ev00__0state >= 6'd25;
wire _guard3426 = ev00__0state <= 6'd25;
wire _guard3427 = _guard3425 & _guard3426;
wire _guard3428 = ev00__0state >= 6'd12;
wire _guard3429 = ev00__0state <= 6'd12;
wire _guard3430 = _guard3428 & _guard3429;
wire _guard3431 = ev00__0state >= 6'd51;
wire _guard3432 = ev00__0state <= 6'd51;
wire _guard3433 = _guard3431 & _guard3432;
wire _guard3434 = ev00__0state >= 6'd38;
wire _guard3435 = ev00__0state <= 6'd38;
wire _guard3436 = _guard3434 & _guard3435;
wire _guard3437 = ev00__0state >= 6'd25;
wire _guard3438 = ev00__0state <= 6'd25;
wire _guard3439 = _guard3437 & _guard3438;
wire _guard3440 = ev00__0state >= 6'd51;
wire _guard3441 = ev00__0state <= 6'd51;
wire _guard3442 = _guard3440 & _guard3441;
wire _guard3443 = ev00__0state >= 6'd12;
wire _guard3444 = ev00__0state <= 6'd12;
wire _guard3445 = _guard3443 & _guard3444;
wire _guard3446 = ev00__0state >= 6'd12;
wire _guard3447 = ev00__0state <= 6'd12;
wire _guard3448 = _guard3446 & _guard3447;
wire _guard3449 = ev00__0state >= 6'd38;
wire _guard3450 = ev00__0state <= 6'd38;
wire _guard3451 = _guard3449 & _guard3450;
wire _guard3452 = ev00__0state >= 6'd25;
wire _guard3453 = ev00__0state <= 6'd25;
wire _guard3454 = _guard3452 & _guard3453;
wire _guard3455 = ev00__0state >= 6'd51;
wire _guard3456 = ev00__0state <= 6'd51;
wire _guard3457 = _guard3455 & _guard3456;
wire _guard3458 = ev00__0state >= 6'd38;
wire _guard3459 = ev00__0state <= 6'd38;
wire _guard3460 = _guard3458 & _guard3459;
wire _guard3461 = ev00__0state >= 6'd25;
wire _guard3462 = ev00__0state <= 6'd25;
wire _guard3463 = _guard3461 & _guard3462;
wire _guard3464 = ev00__0state >= 6'd12;
wire _guard3465 = ev00__0state <= 6'd12;
wire _guard3466 = _guard3464 & _guard3465;
wire _guard3467 = ev00__0state >= 6'd51;
wire _guard3468 = ev00__0state <= 6'd51;
wire _guard3469 = _guard3467 & _guard3468;
wire _guard3470 = ev00__0state >= 6'd12;
wire _guard3471 = ev00__0state <= 6'd12;
wire _guard3472 = _guard3470 & _guard3471;
wire _guard3473 = ev00__0state >= 6'd38;
wire _guard3474 = ev00__0state <= 6'd38;
wire _guard3475 = _guard3473 & _guard3474;
wire _guard3476 = ev00__0state >= 6'd25;
wire _guard3477 = ev00__0state <= 6'd25;
wire _guard3478 = _guard3476 & _guard3477;
wire _guard3479 = ev00__0state >= 6'd51;
wire _guard3480 = ev00__0state <= 6'd51;
wire _guard3481 = _guard3479 & _guard3480;
wire _guard3482 = ev00__0state >= 6'd38;
wire _guard3483 = ev00__0state <= 6'd38;
wire _guard3484 = _guard3482 & _guard3483;
wire _guard3485 = ev00__0state >= 6'd25;
wire _guard3486 = ev00__0state <= 6'd25;
wire _guard3487 = _guard3485 & _guard3486;
wire _guard3488 = ev00__0state >= 6'd12;
wire _guard3489 = ev00__0state <= 6'd12;
wire _guard3490 = _guard3488 & _guard3489;
wire _guard3491 = ev00__0state >= 6'd51;
wire _guard3492 = ev00__0state <= 6'd51;
wire _guard3493 = _guard3491 & _guard3492;
wire _guard3494 = ev00__0state >= 6'd38;
wire _guard3495 = ev00__0state <= 6'd38;
wire _guard3496 = _guard3494 & _guard3495;
wire _guard3497 = ev00__0state >= 6'd12;
wire _guard3498 = ev00__0state <= 6'd12;
wire _guard3499 = _guard3497 & _guard3498;
wire _guard3500 = ev00__0state >= 6'd25;
wire _guard3501 = ev00__0state <= 6'd25;
wire _guard3502 = _guard3500 & _guard3501;
wire _guard3503 = ev00__0state >= 6'd51;
wire _guard3504 = ev00__0state <= 6'd51;
wire _guard3505 = _guard3503 & _guard3504;
wire _guard3506 = ev00__0state >= 6'd51;
wire _guard3507 = ev00__0state <= 6'd51;
wire _guard3508 = _guard3506 & _guard3507;
wire _guard3509 = ev00__0state >= 6'd12;
wire _guard3510 = ev00__0state <= 6'd12;
wire _guard3511 = _guard3509 & _guard3510;
wire _guard3512 = ev00__0state >= 6'd25;
wire _guard3513 = ev00__0state <= 6'd25;
wire _guard3514 = _guard3512 & _guard3513;
wire _guard3515 = ev00__0state >= 6'd38;
wire _guard3516 = ev00__0state <= 6'd38;
wire _guard3517 = _guard3515 & _guard3516;
wire _guard3518 = ev00__0_0;
wire _guard3519 = ev00__0state >= 6'd1;
wire _guard3520 = ev00__0state <= 6'd0;
wire _guard3521 = _guard3519 & _guard3520;
wire _guard3522 = _guard3518 | _guard3521;
wire _guard3523 = ev00__0_0;
wire _guard3524 = ev00__0state >= 6'd1;
wire _guard3525 = ev00__0state <= 6'd0;
wire _guard3526 = _guard3524 & _guard3525;
wire _guard3527 = _guard3523 | _guard3526;
wire _guard3528 = ev00__0_0;
wire _guard3529 = ev00__0state >= 6'd1;
wire _guard3530 = ev00__0state <= 6'd0;
wire _guard3531 = _guard3529 & _guard3530;
wire _guard3532 = _guard3528 | _guard3531;
wire _guard3533 = ev00__0_0;
wire _guard3534 = ev00__0state >= 6'd1;
wire _guard3535 = ev00__0state <= 6'd0;
wire _guard3536 = _guard3534 & _guard3535;
wire _guard3537 = _guard3533 | _guard3536;
wire _guard3538 = ev00__0_0;
wire _guard3539 = ev00__0state >= 6'd1;
wire _guard3540 = ev00__0state <= 6'd0;
wire _guard3541 = _guard3539 & _guard3540;
wire _guard3542 = _guard3538 | _guard3541;
wire _guard3543 = ev00__0state >= 6'd12;
wire _guard3544 = ev00__0state <= 6'd12;
wire _guard3545 = _guard3543 & _guard3544;
wire _guard3546 = ev00__0state >= 6'd26;
wire _guard3547 = ev00__0state <= 6'd26;
wire _guard3548 = _guard3546 & _guard3547;
wire _guard3549 = ev00__0state >= 6'd26;
wire _guard3550 = ev00__0state <= 6'd26;
wire _guard3551 = _guard3549 & _guard3550;
wire _guard3552 = ev00__0state >= 6'd26;
wire _guard3553 = ev00__0state <= 6'd26;
wire _guard3554 = _guard3552 & _guard3553;
wire _guard3555 = ev00__0state >= 6'd26;
wire _guard3556 = ev00__0state <= 6'd26;
wire _guard3557 = _guard3555 & _guard3556;
wire _guard3558 = ev00__0_0;
wire _guard3559 = ev00__0state >= 6'd1;
wire _guard3560 = ev00__0state <= 6'd0;
wire _guard3561 = _guard3559 & _guard3560;
wire _guard3562 = _guard3558 | _guard3561;
wire _guard3563 = ev00__0state >= 6'd7;
wire _guard3564 = ev00__0state <= 6'd7;
wire _guard3565 = _guard3563 & _guard3564;
wire _guard3566 = _guard3562 | _guard3565;
wire _guard3567 = ev00__0state >= 6'd13;
wire _guard3568 = ev00__0state <= 6'd13;
wire _guard3569 = _guard3567 & _guard3568;
wire _guard3570 = _guard3566 | _guard3569;
wire _guard3571 = ev00__0state >= 6'd20;
wire _guard3572 = ev00__0state <= 6'd20;
wire _guard3573 = _guard3571 & _guard3572;
wire _guard3574 = _guard3570 | _guard3573;
wire _guard3575 = ev00__0state >= 6'd26;
wire _guard3576 = ev00__0state <= 6'd26;
wire _guard3577 = _guard3575 & _guard3576;
wire _guard3578 = _guard3574 | _guard3577;
wire _guard3579 = ev00__0state >= 6'd33;
wire _guard3580 = ev00__0state <= 6'd33;
wire _guard3581 = _guard3579 & _guard3580;
wire _guard3582 = _guard3578 | _guard3581;
wire _guard3583 = ev00__0state >= 6'd39;
wire _guard3584 = ev00__0state <= 6'd39;
wire _guard3585 = _guard3583 & _guard3584;
wire _guard3586 = _guard3582 | _guard3585;
wire _guard3587 = ev00__0state >= 6'd46;
wire _guard3588 = ev00__0state <= 6'd46;
wire _guard3589 = _guard3587 & _guard3588;
wire _guard3590 = _guard3586 | _guard3589;
wire _guard3591 = ev00__0state >= 6'd33;
wire _guard3592 = ev00__0state <= 6'd33;
wire _guard3593 = _guard3591 & _guard3592;
wire _guard3594 = ev00__0state >= 6'd39;
wire _guard3595 = ev00__0state <= 6'd39;
wire _guard3596 = _guard3594 & _guard3595;
wire _guard3597 = ev00__0state >= 6'd46;
wire _guard3598 = ev00__0state <= 6'd46;
wire _guard3599 = _guard3597 & _guard3598;
wire _guard3600 = ev00__0state >= 6'd13;
wire _guard3601 = ev00__0state <= 6'd13;
wire _guard3602 = _guard3600 & _guard3601;
wire _guard3603 = ev00__0_0;
wire _guard3604 = ev00__0state >= 6'd1;
wire _guard3605 = ev00__0state <= 6'd0;
wire _guard3606 = _guard3604 & _guard3605;
wire _guard3607 = _guard3603 | _guard3606;
wire _guard3608 = ev00__0state >= 6'd26;
wire _guard3609 = ev00__0state <= 6'd26;
wire _guard3610 = _guard3608 & _guard3609;
wire _guard3611 = ev00__0state >= 6'd7;
wire _guard3612 = ev00__0state <= 6'd7;
wire _guard3613 = _guard3611 & _guard3612;
wire _guard3614 = ev00__0state >= 6'd20;
wire _guard3615 = ev00__0state <= 6'd20;
wire _guard3616 = _guard3614 & _guard3615;
wire _guard3617 = ev00__0state >= 6'd12;
wire _guard3618 = ev00__0state <= 6'd12;
wire _guard3619 = _guard3617 & _guard3618;
wire _guard3620 = ev00__0state >= 6'd39;
wire _guard3621 = ev00__0state <= 6'd39;
wire _guard3622 = _guard3620 & _guard3621;
wire _guard3623 = ev00__0state >= 6'd39;
wire _guard3624 = ev00__0state <= 6'd39;
wire _guard3625 = _guard3623 & _guard3624;
wire _guard3626 = ev00__0state >= 6'd39;
wire _guard3627 = ev00__0state <= 6'd39;
wire _guard3628 = _guard3626 & _guard3627;
wire _guard3629 = ev00__0state >= 6'd39;
wire _guard3630 = ev00__0state <= 6'd39;
wire _guard3631 = _guard3629 & _guard3630;
wire _guard3632 = ev00__0state >= 6'd47;
wire _guard3633 = ev00__0state <= 6'd47;
wire _guard3634 = _guard3632 & _guard3633;
wire _guard3635 = ev00__0state >= 6'd47;
wire _guard3636 = ev00__0state <= 6'd47;
wire _guard3637 = _guard3635 & _guard3636;
wire _guard3638 = ev00__0state >= 6'd47;
wire _guard3639 = ev00__0state <= 6'd47;
wire _guard3640 = _guard3638 & _guard3639;
wire _guard3641 = ev00__0state >= 6'd47;
wire _guard3642 = ev00__0state <= 6'd47;
wire _guard3643 = _guard3641 & _guard3642;
wire _guard3644 = ev00__0state >= 6'd18;
wire _guard3645 = ev00__0state <= 6'd18;
wire _guard3646 = _guard3644 & _guard3645;
wire _guard3647 = ev00__0state >= 6'd51;
wire _guard3648 = ev00__0state <= 6'd51;
wire _guard3649 = _guard3647 & _guard3648;
assign inst44_p4 = inst43_out;
assign inst44_clk = clk;
assign inst44_reset = reset;
assign inst56_p4 = inst43_out;
assign inst56_clk = clk;
assign inst56_reset = reset;
assign inst103_p4 = inst94_out;
assign inst103_clk = clk;
assign inst103_reset = reset;
assign inst138_p6 = inst148_p34;
assign inst138_clk = clk;
assign inst138_p5 = inst148_p33;
assign inst138_p8 = inst148_p36;
assign inst138_reset = reset;
assign inst138_p7 = inst148_p35;
assign inst143_p6 = inst0_p15;
assign inst143_clk = clk;
assign inst143_p5 = inst0_p14;
assign inst143_p8 = inst0_p17;
assign inst143_reset = reset;
assign inst143_p7 = inst0_p16;
assign inst151_p19 = inst2_p48;
assign inst151_p28 = inst2_p57;
assign inst151_p29 = inst2_p58;
assign inst151_p12 = inst2_p41;
assign inst151_p16 = inst2_p45;
assign inst151_p6 = inst2_p35;
assign inst151_p9 = inst2_p38;
assign inst151_p15 = inst2_p44;
assign inst151_p17 = inst2_p46;
assign inst151_p20 = inst2_p49;
assign inst151_p21 = inst2_p50;
assign inst151_p23 = inst2_p52;
assign inst151_clk = clk;
assign inst151_p11 = inst2_p40;
assign inst151_p25 = inst2_p54;
assign inst151_p5 = inst2_p34;
assign inst151_p36 = inst2_p65;
assign inst151_p8 = inst2_p37;
assign inst151_p10 = inst2_p39;
assign inst151_reset = reset;
assign inst151_p7 = inst2_p36;
assign inst151_p13 = inst2_p42;
assign inst151_p18 = inst2_p47;
assign inst151_p30 = inst2_p59;
assign inst151_p24 = inst2_p53;
assign inst151_p32 = inst2_p61;
assign inst151_p14 = inst2_p43;
assign inst151_p26 = inst2_p55;
assign inst151_p31 = inst2_p60;
assign inst151_p27 = inst2_p56;
assign inst151_p33 = inst2_p62;
assign inst151_p22 = inst2_p51;
assign inst151_p34 = inst2_p63;
assign inst151_p35 = inst2_p64;
assign p582 =
  _guard134 ? inst152_p27 :
  32'd0;
assign p573 =
  _guard139 ? inst152_p18 :
  32'd0;
assign p581 =
  _guard144 ? inst152_p26 :
  32'd0;
assign p570 =
  _guard149 ? inst152_p15 :
  32'd0;
assign p572 =
  _guard154 ? inst152_p17 :
  32'd0;
assign p571 =
  _guard159 ? inst152_p16 :
  32'd0;
assign p584 =
  _guard164 ? inst152_p29 :
  32'd0;
assign p585 =
  _guard169 ? inst152_p30 :
  32'd0;
assign p560 =
  _guard174 ? inst152_p5 :
  32'd0;
assign p565 =
  _guard179 ? inst152_p10 :
  32'd0;
assign p574 =
  _guard184 ? inst152_p19 :
  32'd0;
assign p576 =
  _guard189 ? inst152_p21 :
  32'd0;
assign p578 =
  _guard194 ? inst152_p23 :
  32'd0;
assign p562 =
  _guard199 ? inst152_p7 :
  32'd0;
assign p583 =
  _guard204 ? inst152_p28 :
  32'd0;
assign p563 =
  _guard209 ? inst152_p8 :
  32'd0;
assign p566 =
  _guard214 ? inst152_p11 :
  32'd0;
assign p586 =
  _guard219 ? inst152_p31 :
  32'd0;
assign p564 =
  _guard224 ? inst152_p9 :
  32'd0;
assign p567 =
  _guard229 ? inst152_p12 :
  32'd0;
assign p580 =
  _guard234 ? inst152_p25 :
  32'd0;
assign p587 =
  _guard239 ? inst152_p32 :
  32'd0;
assign p577 =
  _guard244 ? inst152_p22 :
  32'd0;
assign p589 =
  _guard249 ? inst152_p34 :
  32'd0;
assign p591 =
  _guard254 ? inst152_p36 :
  32'd0;
assign p561 =
  _guard259 ? inst152_p6 :
  32'd0;
assign p575 =
  _guard264 ? inst152_p20 :
  32'd0;
assign p568 =
  _guard269 ? inst152_p13 :
  32'd0;
assign p579 =
  _guard274 ? inst152_p24 :
  32'd0;
assign p588 =
  _guard279 ? inst152_p33 :
  32'd0;
assign p590 =
  _guard284 ? inst152_p35 :
  32'd0;
assign p569 =
  _guard289 ? inst152_p14 :
  32'd0;
assign inst38_p4 = inst26_out;
assign inst38_clk = clk;
assign inst38_reset = reset;
assign inst41_p6 = inst0_p15;
assign inst41_clk = clk;
assign inst41_p5 = inst0_p14;
assign inst41_p8 = inst0_p17;
assign inst41_reset = reset;
assign inst41_p7 = inst0_p16;
assign inst49_p6 = inst146_p14;
assign inst49_clk = clk;
assign inst49_p5 = inst146_p13;
assign inst49_p8 = inst146_p16;
assign inst49_reset = reset;
assign inst49_p7 = inst146_p15;
assign inst50_p6 = inst0_p15;
assign inst50_clk = clk;
assign inst50_p5 = inst0_p14;
assign inst50_p8 = inst0_p17;
assign inst50_reset = reset;
assign inst50_p7 = inst0_p16;
assign inst71_p6 = inst0_p15;
assign inst71_clk = clk;
assign inst71_p5 = inst0_p14;
assign inst71_p8 = inst0_p17;
assign inst71_reset = reset;
assign inst71_p7 = inst0_p16;
assign inst72_p4 = inst60_out;
assign inst72_clk = clk;
assign inst72_reset = reset;
assign inst74_p6 = inst150_p18;
assign inst74_clk = clk;
assign inst74_p5 = inst150_p17;
assign inst74_p8 = inst150_p20;
assign inst74_reset = reset;
assign inst74_p7 = inst150_p19;
assign inst90_p4 = inst77_out;
assign inst90_clk = clk;
assign inst90_reset = reset;
assign inst117_p6 = inst146_p30;
assign inst117_clk = clk;
assign inst117_p5 = inst146_p29;
assign inst117_p8 = inst146_p32;
assign inst117_reset = reset;
assign inst117_p7 = inst146_p31;
assign inst118_p6 = inst0_p15;
assign inst118_clk = clk;
assign inst118_p5 = inst0_p14;
assign inst118_p8 = inst0_p17;
assign inst118_reset = reset;
assign inst118_p7 = inst0_p16;
assign inst5_p12 = inst1_p27;
assign inst5_p16 = inst1_p31;
assign inst5_p4 = inst1_p19;
assign inst5_p6 = inst1_p21;
assign inst5_p9 = inst1_p24;
assign inst5_p15 = inst1_p30;
assign inst5_p17 = inst1_p32;
assign inst5_clk = clk;
assign inst5_p11 = inst1_p26;
assign inst5_p5 = inst1_p20;
assign inst5_p8 = inst1_p23;
assign inst5_p10 = inst1_p25;
assign inst5_p2 = inst1_p17;
assign inst5_p3 = inst1_p18;
assign inst5_reset = reset;
assign inst5_p7 = inst1_p22;
assign inst5_p13 = inst1_p28;
assign inst5_p14 = inst1_p29;
assign inst21_p4 = inst9_out;
assign inst21_clk = clk;
assign inst21_reset = reset;
assign inst34_p4 = inst26_out;
assign inst34_clk = clk;
assign inst34_reset = reset;
assign inst53_p6 = inst148_p14;
assign inst53_clk = clk;
assign inst53_p5 = inst148_p13;
assign inst53_p8 = inst148_p16;
assign inst53_reset = reset;
assign inst53_p7 = inst148_p15;
assign inst55_p4 = inst43_out;
assign inst55_clk = clk;
assign inst55_reset = reset;
assign inst75_p6 = inst0_p15;
assign inst75_clk = clk;
assign inst75_p5 = inst0_p14;
assign inst75_p8 = inst0_p17;
assign inst75_reset = reset;
assign inst75_p7 = inst0_p16;
assign inst101_p6 = inst0_p15;
assign inst101_clk = clk;
assign inst101_p5 = inst0_p14;
assign inst101_p8 = inst0_p17;
assign inst101_reset = reset;
assign inst101_p7 = inst0_p16;
assign inst140_p4 = inst128_out;
assign inst140_clk = clk;
assign inst140_reset = reset;
assign inst15_p6 = inst146_p6;
assign inst15_clk = clk;
assign inst15_p5 = inst146_p5;
assign inst15_p8 = inst146_p8;
assign inst15_reset = reset;
assign inst15_p7 = inst146_p7;
assign inst16_p6 = inst0_p15;
assign inst16_clk = clk;
assign inst16_p5 = inst0_p14;
assign inst16_p8 = inst0_p17;
assign inst16_reset = reset;
assign inst16_p7 = inst0_p16;
assign inst35_p4 = inst26_out;
assign inst35_clk = clk;
assign inst35_reset = reset;
assign inst61_p4 = inst60_out;
assign inst61_clk = clk;
assign inst61_reset = reset;
assign inst66_p6 = inst146_p18;
assign inst66_clk = clk;
assign inst66_p5 = inst146_p17;
assign inst66_p8 = inst146_p20;
assign inst66_reset = reset;
assign inst66_p7 = inst146_p19;
assign inst85_p4 = inst77_out;
assign inst85_clk = clk;
assign inst85_reset = reset;
assign inst104_p6 = inst148_p26;
assign inst104_clk = clk;
assign inst104_p5 = inst148_p25;
assign inst104_p8 = inst148_p28;
assign inst104_reset = reset;
assign inst104_p7 = inst148_p27;
assign inst137_p4 = inst128_out;
assign inst137_clk = clk;
assign inst137_reset = reset;
assign inst145_p19 = inst2_p48;
assign inst145_p28 = inst2_p57;
assign inst145_p29 = inst2_p58;
assign inst145_p12 = inst2_p41;
assign inst145_p16 = inst2_p45;
assign inst145_p6 = inst2_p35;
assign inst145_p9 = inst2_p38;
assign inst145_p15 = inst2_p44;
assign inst145_p17 = inst2_p46;
assign inst145_p20 = inst2_p49;
assign inst145_p21 = inst2_p50;
assign inst145_p23 = inst2_p52;
assign inst145_clk = clk;
assign inst145_p11 = inst2_p40;
assign inst145_p25 = inst2_p54;
assign inst145_p5 = inst2_p34;
assign inst145_p36 = inst2_p65;
assign inst145_p8 = inst2_p37;
assign inst145_p10 = inst2_p39;
assign inst145_reset = reset;
assign inst145_p7 = inst2_p36;
assign inst145_p13 = inst2_p42;
assign inst145_p18 = inst2_p47;
assign inst145_p30 = inst2_p59;
assign inst145_p24 = inst2_p53;
assign inst145_p32 = inst2_p61;
assign inst145_p14 = inst2_p43;
assign inst145_p26 = inst2_p55;
assign inst145_p31 = inst2_p60;
assign inst145_p27 = inst2_p56;
assign inst145_p33 = inst2_p62;
assign inst145_p22 = inst2_p51;
assign inst145_p34 = inst2_p63;
assign inst145_p35 = inst2_p64;
assign inst8_p12 = inst1_p27;
assign inst8_p16 = inst1_p31;
assign inst8_p4 = inst1_p19;
assign inst8_p6 = inst1_p21;
assign inst8_p9 = inst1_p24;
assign inst8_p15 = inst1_p30;
assign inst8_p17 = inst1_p32;
assign inst8_clk = clk;
assign inst8_p11 = inst1_p26;
assign inst8_p5 = inst1_p20;
assign inst8_p8 = inst1_p23;
assign inst8_p10 = inst1_p25;
assign inst8_p2 = inst1_p17;
assign inst8_p3 = inst1_p18;
assign inst8_reset = reset;
assign inst8_p7 = inst1_p22;
assign inst8_p13 = inst1_p28;
assign inst8_p14 = inst1_p29;
assign inst12_p6 = inst0_p15;
assign inst12_clk = clk;
assign inst12_p5 = inst0_p14;
assign inst12_p8 = inst0_p17;
assign inst12_reset = reset;
assign inst12_p7 = inst0_p16;
assign inst31_p4 = inst26_out;
assign inst31_clk = clk;
assign inst31_reset = reset;
assign inst32_p6 = inst146_p10;
assign inst32_clk = clk;
assign inst32_p5 = inst146_p9;
assign inst32_p8 = inst146_p12;
assign inst32_reset = reset;
assign inst32_p7 = inst146_p11;
assign inst68_p4 = inst60_out;
assign inst68_clk = clk;
assign inst68_reset = reset;
assign inst97_p6 = inst0_p15;
assign inst97_clk = clk;
assign inst97_p5 = inst0_p14;
assign inst97_p8 = inst0_p17;
assign inst97_reset = reset;
assign inst97_p7 = inst0_p16;
assign inst106_p4 = inst94_out;
assign inst106_clk = clk;
assign inst106_reset = reset;
assign inst108_p6 = inst150_p26;
assign inst108_clk = clk;
assign inst108_p5 = inst150_p25;
assign inst108_p8 = inst150_p28;
assign inst108_reset = reset;
assign inst108_p7 = inst150_p27;
assign inst120_p4 = inst111_out;
assign inst120_clk = clk;
assign inst120_reset = reset;
assign inst152_p4 = inst4_out;
assign inst152_clk = clk;
assign inst152_reset = reset;
assign inst3_p19 = p545;
assign inst3_p28 = p554;
assign inst3_p29 = p555;
assign inst3_p12 = p538;
assign inst3_p16 = p542;
assign inst3_p4 = p530;
assign inst3_p6 = p532;
assign inst3_p9 = p535;
assign inst3_p15 = p541;
assign inst3_p17 = p543;
assign inst3_p20 = p546;
assign inst3_p21 = p547;
assign inst3_p23 = p549;
assign inst3_clk = clk;
assign inst3_p11 = p537;
assign inst3_p25 = p551;
assign inst3_p5 = p531;
assign inst3_p8 = p534;
assign inst3_p10 = p536;
assign inst3_p2 = p528;
assign inst3_p3 = p529;
assign inst3_reset = reset;
assign inst3_p7 = p533;
assign inst3_p13 = p539;
assign inst3_p18 = p544;
assign inst3_p30 = p556;
assign inst3_p24 = p550;
assign inst3_p32 = p558;
assign inst3_p14 = p540;
assign inst3_p26 = p552;
assign inst3_p31 = p557;
assign inst3_p27 = p553;
assign inst3_p33 = p559;
assign inst3_p22 = p548;
assign inst25_p4 = inst9_out;
assign inst25_clk = clk;
assign inst25_reset = reset;
assign inst29_p6 = inst0_p15;
assign inst29_clk = clk;
assign inst29_p5 = inst0_p14;
assign inst29_p8 = inst0_p17;
assign inst29_reset = reset;
assign inst29_p7 = inst0_p16;
assign inst43_write_en = _guard1019;
assign inst43_clk = clk;
assign inst43_reset = reset;
assign inst43_in =
  _guard1022 ? inst49_p9 :
  _guard1025 ? inst50_p9 :
  _guard1028 ? inst53_p9 :
  _guard1031 ? inst58_p9 :
  _guard1034 ? inst57_p9 :
  _guard1037 ? inst54_p9 :
  _guard1042 ? inst45_p9 :
  _guard1045 ? inst46_p9 :
  'x;
assign inst94_write_en = _guard1078;
assign inst94_clk = clk;
assign inst94_reset = reset;
assign inst94_in =
  _guard1081 ? inst101_p9 :
  _guard1084 ? inst104_p9 :
  _guard1087 ? inst97_p9 :
  _guard1090 ? inst108_p9 :
  _guard1093 ? inst100_p9 :
  _guard1096 ? inst109_p9 :
  _guard1101 ? inst96_p9 :
  _guard1104 ? inst105_p9 :
  'x;
assign inst95_p4 = inst94_out;
assign inst95_clk = clk;
assign inst95_reset = reset;
assign inst111_write_en = _guard1140;
assign inst111_clk = clk;
assign inst111_reset = reset;
assign inst111_in =
  _guard1143 ? inst117_p9 :
  _guard1146 ? inst118_p9 :
  _guard1149 ? inst125_p9 :
  _guard1152 ? inst114_p9 :
  _guard1155 ? inst126_p9 :
  _guard1158 ? inst121_p9 :
  _guard1163 ? inst113_p9 :
  _guard1166 ? inst122_p9 :
  'x;
assign inst124_p4 = inst111_out;
assign inst124_clk = clk;
assign inst124_reset = reset;
assign inst125_p6 = inst150_p30;
assign inst125_clk = clk;
assign inst125_p5 = inst150_p29;
assign inst125_p8 = inst150_p32;
assign inst125_reset = reset;
assign inst125_p7 = inst150_p31;
assign inst136_p4 = inst128_out;
assign inst136_clk = clk;
assign inst136_reset = reset;
assign inst28_p6 = inst3_p39;
assign inst28_clk = clk;
assign inst28_p5 = inst3_p38;
assign inst28_p8 = inst3_p41;
assign inst28_reset = reset;
assign inst28_p7 = inst3_p40;
assign inst39_p4 = inst26_out;
assign inst39_clk = clk;
assign inst39_reset = reset;
assign inst42_p4 = inst26_out;
assign inst42_clk = clk;
assign inst42_reset = reset;
assign inst51_p4 = inst43_out;
assign inst51_clk = clk;
assign inst51_reset = reset;
assign inst52_p4 = inst43_out;
assign inst52_clk = clk;
assign inst52_reset = reset;
assign inst76_p4 = inst60_out;
assign inst76_clk = clk;
assign inst76_reset = reset;
assign inst82_p4 = inst77_out;
assign inst82_clk = clk;
assign inst82_reset = reset;
assign inst87_p6 = inst148_p22;
assign inst87_clk = clk;
assign inst87_p5 = inst148_p21;
assign inst87_p8 = inst148_p24;
assign inst87_reset = reset;
assign inst87_p7 = inst148_p23;
assign inst116_p4 = inst111_out;
assign inst116_clk = clk;
assign inst116_reset = reset;
assign inst131_p6 = inst0_p15;
assign inst131_clk = clk;
assign inst131_p5 = inst0_p14;
assign inst131_p8 = inst0_p17;
assign inst131_reset = reset;
assign inst131_p7 = inst0_p16;
assign inst132_p4 = inst128_out;
assign inst132_clk = clk;
assign inst132_reset = reset;
assign inst134_p6 = inst146_p34;
assign inst134_clk = clk;
assign inst134_p5 = inst146_p33;
assign inst134_p8 = inst146_p36;
assign inst134_reset = reset;
assign inst134_p7 = inst146_p35;
assign inst139_p6 = inst0_p15;
assign inst139_clk = clk;
assign inst139_p5 = inst0_p14;
assign inst139_p8 = inst0_p17;
assign inst139_reset = reset;
assign inst139_p7 = inst0_p16;
assign inst147_p19 = inst2_p48;
assign inst147_p28 = inst2_p57;
assign inst147_p29 = inst2_p58;
assign inst147_p12 = inst2_p41;
assign inst147_p16 = inst2_p45;
assign inst147_p6 = inst2_p35;
assign inst147_p9 = inst2_p38;
assign inst147_p15 = inst2_p44;
assign inst147_p17 = inst2_p46;
assign inst147_p20 = inst2_p49;
assign inst147_p21 = inst2_p50;
assign inst147_p23 = inst2_p52;
assign inst147_clk = clk;
assign inst147_p11 = inst2_p40;
assign inst147_p25 = inst2_p54;
assign inst147_p5 = inst2_p34;
assign inst147_p36 = inst2_p65;
assign inst147_p8 = inst2_p37;
assign inst147_p10 = inst2_p39;
assign inst147_reset = reset;
assign inst147_p7 = inst2_p36;
assign inst147_p13 = inst2_p42;
assign inst147_p18 = inst2_p47;
assign inst147_p30 = inst2_p59;
assign inst147_p24 = inst2_p53;
assign inst147_p32 = inst2_p61;
assign inst147_p14 = inst2_p43;
assign inst147_p26 = inst2_p55;
assign inst147_p31 = inst2_p60;
assign inst147_p27 = inst2_p56;
assign inst147_p33 = inst2_p62;
assign inst147_p22 = inst2_p51;
assign inst147_p34 = inst2_p63;
assign inst147_p35 = inst2_p64;
assign inst148_p4 = inst4_out;
assign inst148_clk = clk;
assign inst148_reset = reset;
assign inst9_write_en = _guard1408;
assign inst9_clk = clk;
assign inst9_reset = reset;
assign inst9_in =
  _guard1411 ? inst15_p9 :
  _guard1414 ? inst16_p9 :
  _guard1417 ? inst12_p9 :
  _guard1420 ? inst24_p9 :
  _guard1423 ? inst23_p9 :
  _guard1426 ? inst19_p9 :
  _guard1429 ? inst20_p9 :
  _guard1434 ? inst11_p9 :
  'x;
assign inst17_p4 = inst9_out;
assign inst17_clk = clk;
assign inst17_reset = reset;
assign inst48_p4 = inst43_out;
assign inst48_clk = clk;
assign inst48_reset = reset;
assign inst62_p6 = inst3_p47;
assign inst62_clk = clk;
assign inst62_p5 = inst3_p46;
assign inst62_p8 = inst3_p49;
assign inst62_reset = reset;
assign inst62_p7 = inst3_p48;
assign inst70_p6 = inst148_p18;
assign inst70_clk = clk;
assign inst70_p5 = inst148_p17;
assign inst70_p8 = inst148_p20;
assign inst70_reset = reset;
assign inst70_p7 = inst148_p19;
assign inst144_p4 = inst128_out;
assign inst144_clk = clk;
assign inst144_reset = reset;
assign inst150_p4 = inst4_out;
assign inst150_clk = clk;
assign inst150_reset = reset;
assign inst1_clk = clk;
assign inst1_reset = reset;
assign inst24_p6 = inst0_p15;
assign inst24_clk = clk;
assign inst24_p5 = inst0_p14;
assign inst24_p8 = inst0_p17;
assign inst24_reset = reset;
assign inst24_p7 = inst0_p16;
assign inst58_p6 = inst0_p15;
assign inst58_clk = clk;
assign inst58_p5 = inst0_p14;
assign inst58_p8 = inst0_p17;
assign inst58_reset = reset;
assign inst58_p7 = inst0_p16;
assign inst78_p4 = inst77_out;
assign inst78_clk = clk;
assign inst78_reset = reset;
assign inst100_p6 = inst146_p26;
assign inst100_clk = clk;
assign inst100_p5 = inst146_p25;
assign inst100_p8 = inst146_p28;
assign inst100_reset = reset;
assign inst100_p7 = inst146_p27;
assign inst128_write_en = _guard1550;
assign inst128_clk = clk;
assign inst128_reset = reset;
assign inst128_in =
  _guard1553 ? inst138_p9 :
  _guard1556 ? inst143_p9 :
  _guard1559 ? inst131_p9 :
  _guard1562 ? inst134_p9 :
  _guard1565 ? inst139_p9 :
  _guard1570 ? inst130_p9 :
  _guard1573 ? inst135_p9 :
  _guard1576 ? inst142_p9 :
  'x;
assign inst141_p4 = inst128_out;
assign inst141_clk = clk;
assign inst141_reset = reset;
assign inst0_p12 =
  _guard1582 ? inst5_p28 :
  _guard1585 ? inst5_p20 :
  _guard1590 ? inst5_p18 :
  _guard1593 ? inst5_p30 :
  _guard1596 ? inst5_p24 :
  _guard1599 ? inst5_p32 :
  _guard1602 ? inst5_p26 :
  _guard1605 ? inst5_p22 :
  _guard1608 ? inst8_p28 :
  _guard1611 ? inst8_p20 :
  _guard1614 ? inst8_p18 :
  _guard1617 ? inst8_p30 :
  _guard1620 ? inst8_p24 :
  _guard1623 ? inst8_p32 :
  _guard1626 ? inst8_p26 :
  _guard1629 ? inst8_p22 :
  _guard1632 ? inst7_p28 :
  _guard1635 ? inst7_p20 :
  _guard1638 ? inst7_p18 :
  _guard1641 ? inst7_p30 :
  _guard1644 ? inst7_p24 :
  _guard1647 ? inst7_p32 :
  _guard1650 ? inst7_p26 :
  _guard1653 ? inst7_p22 :
  _guard1656 ? inst6_p28 :
  _guard1659 ? inst6_p20 :
  _guard1662 ? inst6_p18 :
  _guard1665 ? inst6_p30 :
  _guard1668 ? inst6_p24 :
  _guard1671 ? inst6_p32 :
  _guard1674 ? inst6_p26 :
  _guard1677 ? inst6_p22 :
  'x;
assign inst0_ev0 = _guard1806;
assign inst0_p9 =
  _guard1809 ? inst44_p6 :
  _guard1812 ? inst56_p6 :
  _guard1815 ? inst103_p6 :
  _guard1818 ? inst90_p6 :
  _guard1821 ? inst35_p6 :
  _guard1824 ? inst61_p6 :
  _guard1827 ? inst137_p6 :
  _guard1830 ? inst31_p6 :
  _guard1833 ? inst120_p6 :
  _guard1836 ? inst95_p6 :
  _guard1839 ? inst124_p6 :
  _guard1842 ? inst39_p6 :
  _guard1845 ? inst52_p6 :
  _guard1848 ? inst82_p6 :
  _guard1851 ? inst116_p6 :
  _guard1854 ? inst48_p6 :
  _guard1857 ? inst78_p6 :
  _guard1860 ? inst141_p6 :
  _guard1863 ? inst27_p6 :
  _guard1866 ? inst65_p6 :
  _guard1869 ? inst133_p6 :
  _guard1872 ? inst129_p6 :
  _guard1875 ? inst73_p6 :
  _guard1878 ? inst69_p6 :
  _guard1881 ? inst107_p6 :
  _guard1884 ? inst112_p6 :
  _guard1887 ? inst14_p6 :
  _guard1890 ? inst18_p6 :
  _guard1893 ? inst22_p6 :
  _guard1896 ? inst86_p6 :
  _guard1901 ? inst10_p6 :
  _guard1904 ? inst99_p6 :
  'x;
assign inst0_clk = clk;
assign inst0_p11 =
  _guard1907 ? inst44_p8 :
  _guard1910 ? inst56_p8 :
  _guard1913 ? inst103_p8 :
  _guard1916 ? inst90_p8 :
  _guard1919 ? inst35_p8 :
  _guard1922 ? inst61_p8 :
  _guard1925 ? inst137_p8 :
  _guard1928 ? inst31_p8 :
  _guard1931 ? inst120_p8 :
  _guard1934 ? inst95_p8 :
  _guard1937 ? inst124_p8 :
  _guard1940 ? inst39_p8 :
  _guard1943 ? inst52_p8 :
  _guard1946 ? inst82_p8 :
  _guard1949 ? inst116_p8 :
  _guard1952 ? inst48_p8 :
  _guard1955 ? inst78_p8 :
  _guard1958 ? inst141_p8 :
  _guard1961 ? inst27_p8 :
  _guard1964 ? inst65_p8 :
  _guard1967 ? inst133_p8 :
  _guard1970 ? inst129_p8 :
  _guard1973 ? inst73_p8 :
  _guard1976 ? inst69_p8 :
  _guard1979 ? inst107_p8 :
  _guard1982 ? inst112_p8 :
  _guard1985 ? inst14_p8 :
  _guard1988 ? inst18_p8 :
  _guard1991 ? inst22_p8 :
  _guard1994 ? inst86_p8 :
  _guard1999 ? inst10_p8 :
  _guard2002 ? inst99_p8 :
  'x;
assign inst0_p8 =
  _guard2005 ? inst44_p5 :
  _guard2008 ? inst56_p5 :
  _guard2011 ? inst103_p5 :
  _guard2014 ? inst90_p5 :
  _guard2017 ? inst35_p5 :
  _guard2020 ? inst61_p5 :
  _guard2023 ? inst137_p5 :
  _guard2026 ? inst31_p5 :
  _guard2029 ? inst120_p5 :
  _guard2032 ? inst95_p5 :
  _guard2035 ? inst124_p5 :
  _guard2038 ? inst39_p5 :
  _guard2041 ? inst52_p5 :
  _guard2044 ? inst82_p5 :
  _guard2047 ? inst116_p5 :
  _guard2050 ? inst48_p5 :
  _guard2053 ? inst78_p5 :
  _guard2056 ? inst141_p5 :
  _guard2059 ? inst27_p5 :
  _guard2062 ? inst65_p5 :
  _guard2065 ? inst133_p5 :
  _guard2068 ? inst129_p5 :
  _guard2071 ? inst73_p5 :
  _guard2074 ? inst69_p5 :
  _guard2077 ? inst107_p5 :
  _guard2080 ? inst112_p5 :
  _guard2083 ? inst14_p5 :
  _guard2086 ? inst18_p5 :
  _guard2089 ? inst22_p5 :
  _guard2092 ? inst86_p5 :
  _guard2097 ? inst10_p5 :
  _guard2100 ? inst99_p5 :
  'x;
assign inst0_p10 =
  _guard2103 ? inst44_p7 :
  _guard2106 ? inst56_p7 :
  _guard2109 ? inst103_p7 :
  _guard2112 ? inst90_p7 :
  _guard2115 ? inst35_p7 :
  _guard2118 ? inst61_p7 :
  _guard2121 ? inst137_p7 :
  _guard2124 ? inst31_p7 :
  _guard2127 ? inst120_p7 :
  _guard2130 ? inst95_p7 :
  _guard2133 ? inst124_p7 :
  _guard2136 ? inst39_p7 :
  _guard2139 ? inst52_p7 :
  _guard2142 ? inst82_p7 :
  _guard2145 ? inst116_p7 :
  _guard2148 ? inst48_p7 :
  _guard2151 ? inst78_p7 :
  _guard2154 ? inst141_p7 :
  _guard2157 ? inst27_p7 :
  _guard2160 ? inst65_p7 :
  _guard2163 ? inst133_p7 :
  _guard2166 ? inst129_p7 :
  _guard2169 ? inst73_p7 :
  _guard2172 ? inst69_p7 :
  _guard2175 ? inst107_p7 :
  _guard2178 ? inst112_p7 :
  _guard2181 ? inst14_p7 :
  _guard2184 ? inst18_p7 :
  _guard2187 ? inst22_p7 :
  _guard2190 ? inst86_p7 :
  _guard2195 ? inst10_p7 :
  _guard2198 ? inst99_p7 :
  'x;
assign inst0_reset = reset;
assign inst0_p13 =
  _guard2203 ? inst5_p19 :
  _guard2206 ? inst5_p29 :
  _guard2209 ? inst5_p21 :
  _guard2212 ? inst5_p23 :
  _guard2215 ? inst5_p25 :
  _guard2218 ? inst5_p31 :
  _guard2221 ? inst5_p27 :
  _guard2224 ? inst5_p33 :
  _guard2227 ? inst8_p19 :
  _guard2230 ? inst8_p29 :
  _guard2233 ? inst8_p21 :
  _guard2236 ? inst8_p23 :
  _guard2239 ? inst8_p25 :
  _guard2242 ? inst8_p31 :
  _guard2245 ? inst8_p27 :
  _guard2248 ? inst8_p33 :
  _guard2251 ? inst7_p19 :
  _guard2254 ? inst7_p29 :
  _guard2257 ? inst7_p21 :
  _guard2260 ? inst7_p23 :
  _guard2263 ? inst7_p25 :
  _guard2266 ? inst7_p31 :
  _guard2269 ? inst7_p27 :
  _guard2272 ? inst7_p33 :
  _guard2275 ? inst6_p19 :
  _guard2278 ? inst6_p29 :
  _guard2281 ? inst6_p21 :
  _guard2284 ? inst6_p23 :
  _guard2287 ? inst6_p25 :
  _guard2290 ? inst6_p31 :
  _guard2293 ? inst6_p27 :
  _guard2296 ? inst6_p33 :
  'x;
assign inst7_p12 = inst1_p27;
assign inst7_p16 = inst1_p31;
assign inst7_p4 = inst1_p19;
assign inst7_p6 = inst1_p21;
assign inst7_p9 = inst1_p24;
assign inst7_p15 = inst1_p30;
assign inst7_p17 = inst1_p32;
assign inst7_clk = clk;
assign inst7_p11 = inst1_p26;
assign inst7_p5 = inst1_p20;
assign inst7_p8 = inst1_p23;
assign inst7_p10 = inst1_p25;
assign inst7_p2 = inst1_p17;
assign inst7_p3 = inst1_p18;
assign inst7_reset = reset;
assign inst7_p7 = inst1_p22;
assign inst7_p13 = inst1_p28;
assign inst7_p14 = inst1_p29;
assign inst23_p6 = inst150_p6;
assign inst23_clk = clk;
assign inst23_p5 = inst150_p5;
assign inst23_p8 = inst150_p8;
assign inst23_reset = reset;
assign inst23_p7 = inst150_p7;
assign inst27_p4 = inst26_out;
assign inst27_clk = clk;
assign inst27_reset = reset;
assign inst30_p4 = inst26_out;
assign inst30_clk = clk;
assign inst30_reset = reset;
assign inst57_p6 = inst150_p14;
assign inst57_clk = clk;
assign inst57_p5 = inst150_p13;
assign inst57_p8 = inst150_p16;
assign inst57_reset = reset;
assign inst57_p7 = inst150_p15;
assign inst59_p4 = inst43_out;
assign inst59_clk = clk;
assign inst59_reset = reset;
assign inst65_p4 = inst60_out;
assign inst65_clk = clk;
assign inst65_reset = reset;
assign inst80_p6 = inst0_p15;
assign inst80_clk = clk;
assign inst80_p5 = inst0_p14;
assign inst80_p8 = inst0_p17;
assign inst80_reset = reset;
assign inst80_p7 = inst0_p16;
assign inst114_p6 = inst0_p15;
assign inst114_clk = clk;
assign inst114_p5 = inst0_p14;
assign inst114_p8 = inst0_p17;
assign inst114_reset = reset;
assign inst114_p7 = inst0_p16;
assign inst126_p6 = inst0_p15;
assign inst126_clk = clk;
assign inst126_p5 = inst0_p14;
assign inst126_p8 = inst0_p17;
assign inst126_reset = reset;
assign inst126_p7 = inst0_p16;
assign inst130_p6 = inst3_p63;
assign inst130_clk = clk;
assign inst130_p5 = inst3_p62;
assign inst130_p8 = inst3_p65;
assign inst130_reset = reset;
assign inst130_p7 = inst3_p64;
assign inst133_p4 = inst128_out;
assign inst133_clk = clk;
assign inst133_reset = reset;
assign inst135_p6 = inst0_p15;
assign inst135_clk = clk;
assign inst135_p5 = inst0_p14;
assign inst135_p8 = inst0_p17;
assign inst135_reset = reset;
assign inst135_p7 = inst0_p16;
assign inst142_p6 = inst150_p34;
assign inst142_clk = clk;
assign inst142_p5 = inst150_p33;
assign inst142_p8 = inst150_p36;
assign inst142_reset = reset;
assign inst142_p7 = inst150_p35;
assign inst146_p4 = inst4_out;
assign inst146_clk = clk;
assign inst146_reset = reset;
assign inst19_p6 = inst148_p6;
assign inst19_clk = clk;
assign inst19_p5 = inst148_p5;
assign inst19_p8 = inst148_p8;
assign inst19_reset = reset;
assign inst19_p7 = inst148_p7;
assign inst40_p6 = inst150_p10;
assign inst40_clk = clk;
assign inst40_p5 = inst150_p9;
assign inst40_p8 = inst150_p12;
assign inst40_reset = reset;
assign inst40_p7 = inst150_p11;
assign inst64_p4 = inst60_out;
assign inst64_clk = clk;
assign inst64_reset = reset;
assign inst83_p6 = inst146_p22;
assign inst83_clk = clk;
assign inst83_p5 = inst146_p21;
assign inst83_p8 = inst146_p24;
assign inst83_reset = reset;
assign inst83_p7 = inst146_p23;
assign inst109_p6 = inst0_p15;
assign inst109_clk = clk;
assign inst109_p5 = inst0_p14;
assign inst109_p8 = inst0_p17;
assign inst109_reset = reset;
assign inst109_p7 = inst0_p16;
assign inst129_p4 = inst128_out;
assign inst129_clk = clk;
assign inst129_reset = reset;
assign ev00_clk = clk;
assign ev00_go = ev0;
assign ev00_reset = reset;
assign inst54_p6 = inst0_p15;
assign inst54_clk = clk;
assign inst54_p5 = inst0_p14;
assign inst54_p8 = inst0_p17;
assign inst54_reset = reset;
assign inst54_p7 = inst0_p16;
assign inst73_p4 = inst60_out;
assign inst73_clk = clk;
assign inst73_reset = reset;
assign inst88_p6 = inst0_p15;
assign inst88_clk = clk;
assign inst88_p5 = inst0_p14;
assign inst88_p8 = inst0_p17;
assign inst88_reset = reset;
assign inst88_p7 = inst0_p16;
assign inst98_p4 = inst94_out;
assign inst98_clk = clk;
assign inst98_reset = reset;
assign inst102_p4 = inst94_out;
assign inst102_clk = clk;
assign inst102_reset = reset;
assign inst45_p6 = inst3_p43;
assign inst45_clk = clk;
assign inst45_p5 = inst3_p42;
assign inst45_p8 = inst3_p45;
assign inst45_reset = reset;
assign inst45_p7 = inst3_p44;
assign inst46_p6 = inst0_p15;
assign inst46_clk = clk;
assign inst46_p5 = inst0_p14;
assign inst46_p8 = inst0_p17;
assign inst46_reset = reset;
assign inst46_p7 = inst0_p16;
assign inst47_p4 = inst43_out;
assign inst47_clk = clk;
assign inst47_reset = reset;
assign inst69_p4 = inst60_out;
assign inst69_clk = clk;
assign inst69_reset = reset;
assign inst84_p6 = inst0_p15;
assign inst84_clk = clk;
assign inst84_p5 = inst0_p14;
assign inst84_p8 = inst0_p17;
assign inst84_reset = reset;
assign inst84_p7 = inst0_p16;
assign inst96_p6 = inst3_p55;
assign inst96_clk = clk;
assign inst96_p5 = inst3_p54;
assign inst96_p8 = inst3_p57;
assign inst96_reset = reset;
assign inst96_p7 = inst3_p56;
assign inst107_p4 = inst94_out;
assign inst107_clk = clk;
assign inst107_reset = reset;
assign inst112_p4 = inst111_out;
assign inst112_clk = clk;
assign inst112_reset = reset;
assign inst6_p12 = inst1_p27;
assign inst6_p16 = inst1_p31;
assign inst6_p4 = inst1_p19;
assign inst6_p6 = inst1_p21;
assign inst6_p9 = inst1_p24;
assign inst6_p15 = inst1_p30;
assign inst6_p17 = inst1_p32;
assign inst6_clk = clk;
assign inst6_p11 = inst1_p26;
assign inst6_p5 = inst1_p20;
assign inst6_p8 = inst1_p23;
assign inst6_p10 = inst1_p25;
assign inst6_p2 = inst1_p17;
assign inst6_p3 = inst1_p18;
assign inst6_reset = reset;
assign inst6_p7 = inst1_p22;
assign inst6_p13 = inst1_p28;
assign inst6_p14 = inst1_p29;
assign inst20_p6 = inst0_p15;
assign inst20_clk = clk;
assign inst20_p5 = inst0_p14;
assign inst20_p8 = inst0_p17;
assign inst20_reset = reset;
assign inst20_p7 = inst0_p16;
assign inst33_p6 = inst0_p15;
assign inst33_clk = clk;
assign inst33_p5 = inst0_p14;
assign inst33_p8 = inst0_p17;
assign inst33_reset = reset;
assign inst33_p7 = inst0_p16;
assign inst77_write_en = _guard2798;
assign inst77_clk = clk;
assign inst77_reset = reset;
assign inst77_in =
  _guard2801 ? inst87_p9 :
  _guard2804 ? inst80_p9 :
  _guard2807 ? inst83_p9 :
  _guard2810 ? inst88_p9 :
  _guard2813 ? inst84_p9 :
  _guard2818 ? inst79_p9 :
  _guard2821 ? inst91_p9 :
  _guard2824 ? inst92_p9 :
  'x;
assign inst79_p6 = inst3_p51;
assign inst79_clk = clk;
assign inst79_p5 = inst3_p50;
assign inst79_p8 = inst3_p53;
assign inst79_reset = reset;
assign inst79_p7 = inst3_p52;
assign inst93_p4 = inst77_out;
assign inst93_clk = clk;
assign inst93_reset = reset;
assign inst115_p4 = inst111_out;
assign inst115_clk = clk;
assign inst115_reset = reset;
assign inst121_p6 = inst148_p30;
assign inst121_clk = clk;
assign inst121_p5 = inst148_p29;
assign inst121_p8 = inst148_p32;
assign inst121_reset = reset;
assign inst121_p7 = inst148_p31;
assign inst123_p4 = inst111_out;
assign inst123_clk = clk;
assign inst123_reset = reset;
assign inst149_p19 = inst2_p48;
assign inst149_p28 = inst2_p57;
assign inst149_p29 = inst2_p58;
assign inst149_p12 = inst2_p41;
assign inst149_p16 = inst2_p45;
assign inst149_p6 = inst2_p35;
assign inst149_p9 = inst2_p38;
assign inst149_p15 = inst2_p44;
assign inst149_p17 = inst2_p46;
assign inst149_p20 = inst2_p49;
assign inst149_p21 = inst2_p50;
assign inst149_p23 = inst2_p52;
assign inst149_clk = clk;
assign inst149_p11 = inst2_p40;
assign inst149_p25 = inst2_p54;
assign inst149_p5 = inst2_p34;
assign inst149_p36 = inst2_p65;
assign inst149_p8 = inst2_p37;
assign inst149_p10 = inst2_p39;
assign inst149_reset = reset;
assign inst149_p7 = inst2_p36;
assign inst149_p13 = inst2_p42;
assign inst149_p18 = inst2_p47;
assign inst149_p30 = inst2_p59;
assign inst149_p24 = inst2_p53;
assign inst149_p32 = inst2_p61;
assign inst149_p14 = inst2_p43;
assign inst149_p26 = inst2_p55;
assign inst149_p31 = inst2_p60;
assign inst149_p27 = inst2_p56;
assign inst149_p33 = inst2_p62;
assign inst149_p22 = inst2_p51;
assign inst149_p34 = inst2_p63;
assign inst149_p35 = inst2_p64;
assign inst14_p4 = inst9_out;
assign inst14_clk = clk;
assign inst14_reset = reset;
assign inst18_p4 = inst9_out;
assign inst18_clk = clk;
assign inst18_reset = reset;
assign inst22_p4 = inst9_out;
assign inst22_clk = clk;
assign inst22_reset = reset;
assign inst26_write_en = _guard3003;
assign inst26_clk = clk;
assign inst26_reset = reset;
assign inst26_in =
  _guard3006 ? inst41_p9 :
  _guard3009 ? inst32_p9 :
  _guard3012 ? inst29_p9 :
  _guard3017 ? inst28_p9 :
  _guard3020 ? inst40_p9 :
  _guard3023 ? inst33_p9 :
  _guard3026 ? inst37_p9 :
  _guard3029 ? inst36_p9 :
  'x;
assign inst37_p6 = inst0_p15;
assign inst37_clk = clk;
assign inst37_p5 = inst0_p14;
assign inst37_p8 = inst0_p17;
assign inst37_reset = reset;
assign inst37_p7 = inst0_p16;
assign inst63_p6 = inst0_p15;
assign inst63_clk = clk;
assign inst63_p5 = inst0_p14;
assign inst63_p8 = inst0_p17;
assign inst63_reset = reset;
assign inst63_p7 = inst0_p16;
assign inst67_p6 = inst0_p15;
assign inst67_clk = clk;
assign inst67_p5 = inst0_p14;
assign inst67_p8 = inst0_p17;
assign inst67_reset = reset;
assign inst67_p7 = inst0_p16;
assign inst86_p4 = inst77_out;
assign inst86_clk = clk;
assign inst86_reset = reset;
assign inst89_p4 = inst77_out;
assign inst89_clk = clk;
assign inst89_reset = reset;
assign inst105_p6 = inst0_p15;
assign inst105_clk = clk;
assign inst105_p5 = inst0_p14;
assign inst105_p8 = inst0_p17;
assign inst105_reset = reset;
assign inst105_p7 = inst0_p16;
assign inst113_p6 = inst3_p59;
assign inst113_clk = clk;
assign inst113_p5 = inst3_p58;
assign inst113_p8 = inst3_p61;
assign inst113_reset = reset;
assign inst113_p7 = inst3_p60;
assign inst119_p4 = inst111_out;
assign inst119_clk = clk;
assign inst119_reset = reset;
assign inst122_p6 = inst0_p15;
assign inst122_clk = clk;
assign inst122_p5 = inst0_p14;
assign inst122_p8 = inst0_p17;
assign inst122_reset = reset;
assign inst122_p7 = inst0_p16;
assign inst127_p4 = inst111_out;
assign inst127_clk = clk;
assign inst127_reset = reset;
assign inst2_p19 =
  _guard3124 ? inst85_p6 :
  _guard3127 ? inst93_p6 :
  _guard3130 ? inst89_p6 :
  _guard3133 ? inst81_p6 :
  'x;
assign inst2_p28 =
  _guard3136 ? inst115_p7 :
  _guard3139 ? inst123_p7 :
  _guard3142 ? inst119_p7 :
  _guard3145 ? inst127_p7 :
  'x;
assign inst2_p29 =
  _guard3148 ? inst115_p8 :
  _guard3151 ? inst123_p8 :
  _guard3154 ? inst119_p8 :
  _guard3157 ? inst127_p8 :
  'x;
assign inst2_p12 =
  _guard3160 ? inst55_p7 :
  _guard3163 ? inst51_p7 :
  _guard3166 ? inst59_p7 :
  _guard3169 ? inst47_p7 :
  'x;
assign inst2_p16 =
  _guard3172 ? inst72_p7 :
  _guard3175 ? inst68_p7 :
  _guard3178 ? inst76_p7 :
  _guard3181 ? inst64_p7 :
  'x;
assign inst2_p4 =
  _guard3184 ? inst21_p7 :
  _guard3187 ? inst25_p7 :
  _guard3190 ? inst17_p7 :
  _guard3193 ? inst13_p7 :
  'x;
assign inst2_p6 =
  _guard3196 ? inst38_p5 :
  _guard3199 ? inst34_p5 :
  _guard3202 ? inst42_p5 :
  _guard3205 ? inst30_p5 :
  'x;
assign inst2_p9 =
  _guard3208 ? inst38_p8 :
  _guard3211 ? inst34_p8 :
  _guard3214 ? inst42_p8 :
  _guard3217 ? inst30_p8 :
  'x;
assign inst2_p15 =
  _guard3220 ? inst72_p6 :
  _guard3223 ? inst68_p6 :
  _guard3226 ? inst76_p6 :
  _guard3229 ? inst64_p6 :
  'x;
assign inst2_p17 =
  _guard3232 ? inst72_p8 :
  _guard3235 ? inst68_p8 :
  _guard3238 ? inst76_p8 :
  _guard3241 ? inst64_p8 :
  'x;
assign inst2_p20 =
  _guard3244 ? inst85_p7 :
  _guard3247 ? inst93_p7 :
  _guard3250 ? inst89_p7 :
  _guard3253 ? inst81_p7 :
  'x;
assign inst2_p21 =
  _guard3256 ? inst85_p8 :
  _guard3259 ? inst93_p8 :
  _guard3262 ? inst89_p8 :
  _guard3265 ? inst81_p8 :
  'x;
assign inst2_p23 =
  _guard3268 ? inst106_p6 :
  _guard3271 ? inst98_p6 :
  _guard3274 ? inst102_p6 :
  _guard3277 ? inst110_p6 :
  'x;
assign inst2_clk = clk;
assign inst2_p11 =
  _guard3280 ? inst55_p6 :
  _guard3283 ? inst51_p6 :
  _guard3286 ? inst59_p6 :
  _guard3289 ? inst47_p6 :
  'x;
assign inst2_p25 =
  _guard3292 ? inst106_p8 :
  _guard3295 ? inst98_p8 :
  _guard3298 ? inst102_p8 :
  _guard3301 ? inst110_p8 :
  'x;
assign inst2_p5 =
  _guard3304 ? inst21_p8 :
  _guard3307 ? inst25_p8 :
  _guard3310 ? inst17_p8 :
  _guard3313 ? inst13_p8 :
  'x;
assign inst2_p8 =
  _guard3316 ? inst38_p7 :
  _guard3319 ? inst34_p7 :
  _guard3322 ? inst42_p7 :
  _guard3325 ? inst30_p7 :
  'x;
assign inst2_p10 =
  _guard3328 ? inst55_p5 :
  _guard3331 ? inst51_p5 :
  _guard3334 ? inst59_p5 :
  _guard3337 ? inst47_p5 :
  'x;
assign inst2_p2 =
  _guard3340 ? inst21_p5 :
  _guard3343 ? inst25_p5 :
  _guard3346 ? inst17_p5 :
  _guard3349 ? inst13_p5 :
  'x;
assign inst2_p3 =
  _guard3352 ? inst21_p6 :
  _guard3355 ? inst25_p6 :
  _guard3358 ? inst17_p6 :
  _guard3361 ? inst13_p6 :
  'x;
assign inst2_reset = reset;
assign inst2_p7 =
  _guard3364 ? inst38_p6 :
  _guard3367 ? inst34_p6 :
  _guard3370 ? inst42_p6 :
  _guard3373 ? inst30_p6 :
  'x;
assign inst2_p13 =
  _guard3376 ? inst55_p8 :
  _guard3379 ? inst51_p8 :
  _guard3382 ? inst59_p8 :
  _guard3385 ? inst47_p8 :
  'x;
assign inst2_p18 =
  _guard3388 ? inst85_p5 :
  _guard3391 ? inst93_p5 :
  _guard3394 ? inst89_p5 :
  _guard3397 ? inst81_p5 :
  'x;
assign inst2_p30 =
  _guard3400 ? inst140_p5 :
  _guard3403 ? inst136_p5 :
  _guard3406 ? inst132_p5 :
  _guard3409 ? inst144_p5 :
  'x;
assign inst2_p24 =
  _guard3412 ? inst106_p7 :
  _guard3415 ? inst98_p7 :
  _guard3418 ? inst102_p7 :
  _guard3421 ? inst110_p7 :
  'x;
assign inst2_p32 =
  _guard3424 ? inst140_p7 :
  _guard3427 ? inst136_p7 :
  _guard3430 ? inst132_p7 :
  _guard3433 ? inst144_p7 :
  'x;
assign inst2_p14 =
  _guard3436 ? inst72_p5 :
  _guard3439 ? inst68_p5 :
  _guard3442 ? inst76_p5 :
  _guard3445 ? inst64_p5 :
  'x;
assign inst2_p26 =
  _guard3448 ? inst115_p5 :
  _guard3451 ? inst123_p5 :
  _guard3454 ? inst119_p5 :
  _guard3457 ? inst127_p5 :
  'x;
assign inst2_p31 =
  _guard3460 ? inst140_p6 :
  _guard3463 ? inst136_p6 :
  _guard3466 ? inst132_p6 :
  _guard3469 ? inst144_p6 :
  'x;
assign inst2_p27 =
  _guard3472 ? inst115_p6 :
  _guard3475 ? inst123_p6 :
  _guard3478 ? inst119_p6 :
  _guard3481 ? inst127_p6 :
  'x;
assign inst2_p33 =
  _guard3484 ? inst140_p8 :
  _guard3487 ? inst136_p8 :
  _guard3490 ? inst132_p8 :
  _guard3493 ? inst144_p8 :
  'x;
assign inst2_p22 =
  _guard3496 ? inst106_p5 :
  _guard3499 ? inst98_p5 :
  _guard3502 ? inst102_p5 :
  _guard3505 ? inst110_p5 :
  'x;
assign inst4_clk = clk;
assign inst4_reset = reset;
assign inst4_in =
  _guard3508 ? inst151_p37 :
  _guard3511 ? inst145_p37 :
  _guard3514 ? inst147_p37 :
  _guard3517 ? inst149_p37 :
  'x;
assign inst10_p4 = inst9_out;
assign inst10_clk = clk;
assign inst10_reset = reset;
assign inst11_p6 = inst3_p35;
assign inst11_clk = clk;
assign inst11_p5 = inst3_p34;
assign inst11_p8 = inst3_p37;
assign inst11_reset = reset;
assign inst11_p7 = inst3_p36;
assign inst13_p4 = inst9_out;
assign inst13_clk = clk;
assign inst13_reset = reset;
assign inst36_p6 = inst148_p10;
assign inst36_clk = clk;
assign inst36_p5 = inst148_p9;
assign inst36_p8 = inst148_p12;
assign inst36_reset = reset;
assign inst36_p7 = inst148_p11;
assign inst60_write_en = _guard3590;
assign inst60_clk = clk;
assign inst60_reset = reset;
assign inst60_in =
  _guard3593 ? inst71_p9 :
  _guard3596 ? inst74_p9 :
  _guard3599 ? inst75_p9 :
  _guard3602 ? inst66_p9 :
  _guard3607 ? inst62_p9 :
  _guard3610 ? inst70_p9 :
  _guard3613 ? inst63_p9 :
  _guard3616 ? inst67_p9 :
  'x;
assign inst81_p4 = inst77_out;
assign inst81_clk = clk;
assign inst81_reset = reset;
assign inst91_p6 = inst150_p22;
assign inst91_clk = clk;
assign inst91_p5 = inst150_p21;
assign inst91_p8 = inst150_p24;
assign inst91_reset = reset;
assign inst91_p7 = inst150_p23;
assign inst92_p6 = inst0_p15;
assign inst92_clk = clk;
assign inst92_p5 = inst0_p14;
assign inst92_p8 = inst0_p17;
assign inst92_reset = reset;
assign inst92_p7 = inst0_p16;
assign inst99_p4 = inst94_out;
assign inst99_clk = clk;
assign inst99_reset = reset;
assign inst110_p4 = inst94_out;
assign inst110_clk = clk;
assign inst110_reset = reset;
// COMPONENT END: comp94
endmodule
module comp95(
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  input logic [31:0] p37,
  input logic [31:0] p38,
  input logic [31:0] p39,
  output logic [1023:0] p40,
  input logic ev0,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp95
logic [5:0] ev00__0state;
logic ev00__0_0;
logic [5:0] ev00__1state;
logic ev00__1_0;
logic ev00_clk;
logic ev00_reset;
logic ev00_go;
logic ev00_done;
logic [31:0] inst0_p528;
logic [31:0] inst0_p529;
logic [31:0] inst0_p530;
logic [31:0] inst0_p531;
logic [31:0] inst0_p532;
logic [31:0] inst0_p533;
logic [31:0] inst0_p534;
logic [31:0] inst0_p535;
logic [31:0] inst0_p536;
logic [31:0] inst0_p537;
logic [31:0] inst0_p538;
logic [31:0] inst0_p539;
logic [31:0] inst0_p540;
logic [31:0] inst0_p541;
logic [31:0] inst0_p542;
logic [31:0] inst0_p543;
logic [31:0] inst0_p544;
logic [31:0] inst0_p545;
logic [31:0] inst0_p546;
logic [31:0] inst0_p547;
logic [31:0] inst0_p548;
logic [31:0] inst0_p549;
logic [31:0] inst0_p550;
logic [31:0] inst0_p551;
logic [31:0] inst0_p552;
logic [31:0] inst0_p553;
logic [31:0] inst0_p554;
logic [31:0] inst0_p555;
logic [31:0] inst0_p556;
logic [31:0] inst0_p557;
logic [31:0] inst0_p558;
logic [31:0] inst0_p559;
logic [31:0] inst0_p560;
logic [31:0] inst0_p561;
logic [31:0] inst0_p562;
logic [31:0] inst0_p563;
logic [31:0] inst0_p564;
logic [31:0] inst0_p565;
logic [31:0] inst0_p566;
logic [31:0] inst0_p567;
logic [31:0] inst0_p568;
logic [31:0] inst0_p569;
logic [31:0] inst0_p570;
logic [31:0] inst0_p571;
logic [31:0] inst0_p572;
logic [31:0] inst0_p573;
logic [31:0] inst0_p574;
logic [31:0] inst0_p575;
logic [31:0] inst0_p576;
logic [31:0] inst0_p577;
logic [31:0] inst0_p578;
logic [31:0] inst0_p579;
logic [31:0] inst0_p580;
logic [31:0] inst0_p581;
logic [31:0] inst0_p582;
logic [31:0] inst0_p583;
logic [31:0] inst0_p584;
logic [31:0] inst0_p585;
logic [31:0] inst0_p586;
logic [31:0] inst0_p587;
logic [31:0] inst0_p588;
logic [31:0] inst0_p589;
logic [31:0] inst0_p590;
logic [31:0] inst0_p591;
logic inst0_ev0;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_p7;
logic [31:0] inst1_p8;
logic [31:0] inst1_p9;
logic [31:0] inst1_p10;
logic [31:0] inst1_p11;
logic [31:0] inst1_p12;
logic [31:0] inst1_p13;
logic [31:0] inst1_p14;
logic [31:0] inst1_p15;
logic [31:0] inst1_p16;
logic [31:0] inst1_p17;
logic [31:0] inst1_p18;
logic [31:0] inst1_p19;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic [31:0] inst1_p30;
logic [31:0] inst1_p31;
logic [31:0] inst1_p32;
logic [31:0] inst1_p33;
logic [31:0] inst1_p34;
logic [31:0] inst1_p35;
logic [31:0] inst1_p36;
logic [31:0] inst1_p37;
logic [31:0] inst1_p38;
logic [1023:0] inst1_p39;
logic inst1_clk;
logic inst1_reset;
counter_chain_2_52 ev00 (
    ._0_0(ev00__0_0),
    ._0state(ev00__0state),
    ._1_0(ev00__1_0),
    ._1state(ev00__1state),
    .clk(ev00_clk),
    .done(ev00_done),
    .go(ev00_go),
    .reset(ev00_reset)
);
comp94 inst0 (
    .clk(inst0_clk),
    .ev0(inst0_ev0),
    .p528(inst0_p528),
    .p529(inst0_p529),
    .p530(inst0_p530),
    .p531(inst0_p531),
    .p532(inst0_p532),
    .p533(inst0_p533),
    .p534(inst0_p534),
    .p535(inst0_p535),
    .p536(inst0_p536),
    .p537(inst0_p537),
    .p538(inst0_p538),
    .p539(inst0_p539),
    .p540(inst0_p540),
    .p541(inst0_p541),
    .p542(inst0_p542),
    .p543(inst0_p543),
    .p544(inst0_p544),
    .p545(inst0_p545),
    .p546(inst0_p546),
    .p547(inst0_p547),
    .p548(inst0_p548),
    .p549(inst0_p549),
    .p550(inst0_p550),
    .p551(inst0_p551),
    .p552(inst0_p552),
    .p553(inst0_p553),
    .p554(inst0_p554),
    .p555(inst0_p555),
    .p556(inst0_p556),
    .p557(inst0_p557),
    .p558(inst0_p558),
    .p559(inst0_p559),
    .p560(inst0_p560),
    .p561(inst0_p561),
    .p562(inst0_p562),
    .p563(inst0_p563),
    .p564(inst0_p564),
    .p565(inst0_p565),
    .p566(inst0_p566),
    .p567(inst0_p567),
    .p568(inst0_p568),
    .p569(inst0_p569),
    .p570(inst0_p570),
    .p571(inst0_p571),
    .p572(inst0_p572),
    .p573(inst0_p573),
    .p574(inst0_p574),
    .p575(inst0_p575),
    .p576(inst0_p576),
    .p577(inst0_p577),
    .p578(inst0_p578),
    .p579(inst0_p579),
    .p580(inst0_p580),
    .p581(inst0_p581),
    .p582(inst0_p582),
    .p583(inst0_p583),
    .p584(inst0_p584),
    .p585(inst0_p585),
    .p586(inst0_p586),
    .p587(inst0_p587),
    .p588(inst0_p588),
    .p589(inst0_p589),
    .p590(inst0_p590),
    .p591(inst0_p591),
    .reset(inst0_reset)
);
comp91 inst1 (
    .clk(inst1_clk),
    .p10(inst1_p10),
    .p11(inst1_p11),
    .p12(inst1_p12),
    .p13(inst1_p13),
    .p14(inst1_p14),
    .p15(inst1_p15),
    .p16(inst1_p16),
    .p17(inst1_p17),
    .p18(inst1_p18),
    .p19(inst1_p19),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .p30(inst1_p30),
    .p31(inst1_p31),
    .p32(inst1_p32),
    .p33(inst1_p33),
    .p34(inst1_p34),
    .p35(inst1_p35),
    .p36(inst1_p36),
    .p37(inst1_p37),
    .p38(inst1_p38),
    .p39(inst1_p39),
    .p7(inst1_p7),
    .p8(inst1_p8),
    .p9(inst1_p9),
    .reset(inst1_reset)
);
wire _guard0 = 1;
wire _guard1 = ev00__1_0;
wire _guard2 = ev00__1state >= 6'd1;
wire _guard3 = ev00__1state <= 6'd0;
wire _guard4 = _guard2 & _guard3;
wire _guard5 = _guard1 | _guard4;
wire _guard6 = ev00__1_0;
wire _guard7 = ev00__1state >= 6'd1;
wire _guard8 = ev00__1state <= 6'd0;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = _guard6 | _guard9;
wire _guard11 = ev00__1_0;
wire _guard12 = ev00__1state >= 6'd1;
wire _guard13 = ev00__1state <= 6'd0;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = _guard11 | _guard14;
wire _guard16 = ev00__1_0;
wire _guard17 = ev00__1state >= 6'd1;
wire _guard18 = ev00__1state <= 6'd0;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = _guard16 | _guard19;
wire _guard21 = ev00__1_0;
wire _guard22 = ev00__1state >= 6'd1;
wire _guard23 = ev00__1state <= 6'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard21 | _guard24;
wire _guard26 = ev00__1_0;
wire _guard27 = ev00__1state >= 6'd1;
wire _guard28 = ev00__1state <= 6'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard26 | _guard29;
wire _guard31 = ev00__1_0;
wire _guard32 = ev00__1state >= 6'd1;
wire _guard33 = ev00__1state <= 6'd0;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = _guard31 | _guard34;
wire _guard36 = ev00__1_0;
wire _guard37 = ev00__1state >= 6'd1;
wire _guard38 = ev00__1state <= 6'd0;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = _guard36 | _guard39;
wire _guard41 = ev00__1_0;
wire _guard42 = ev00__1state >= 6'd1;
wire _guard43 = ev00__1state <= 6'd0;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = _guard41 | _guard44;
wire _guard46 = ev00__1_0;
wire _guard47 = ev00__1state >= 6'd1;
wire _guard48 = ev00__1state <= 6'd0;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = _guard46 | _guard49;
wire _guard51 = ev00__1_0;
wire _guard52 = ev00__1state >= 6'd1;
wire _guard53 = ev00__1state <= 6'd0;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = _guard51 | _guard54;
wire _guard56 = ev00__1_0;
wire _guard57 = ev00__1state >= 6'd1;
wire _guard58 = ev00__1state <= 6'd0;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = _guard56 | _guard59;
wire _guard61 = ev00__1_0;
wire _guard62 = ev00__1state >= 6'd1;
wire _guard63 = ev00__1state <= 6'd0;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = _guard61 | _guard64;
wire _guard66 = ev00__1_0;
wire _guard67 = ev00__1state >= 6'd1;
wire _guard68 = ev00__1state <= 6'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = _guard66 | _guard69;
wire _guard71 = ev00__1_0;
wire _guard72 = ev00__1state >= 6'd1;
wire _guard73 = ev00__1state <= 6'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard71 | _guard74;
wire _guard76 = ev00__1_0;
wire _guard77 = ev00__1state >= 6'd1;
wire _guard78 = ev00__1state <= 6'd0;
wire _guard79 = _guard77 & _guard78;
wire _guard80 = _guard76 | _guard79;
wire _guard81 = ev00__1_0;
wire _guard82 = ev00__1state >= 6'd1;
wire _guard83 = ev00__1state <= 6'd0;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = _guard81 | _guard84;
wire _guard86 = ev00__1_0;
wire _guard87 = ev00__1state >= 6'd1;
wire _guard88 = ev00__1state <= 6'd0;
wire _guard89 = _guard87 & _guard88;
wire _guard90 = _guard86 | _guard89;
wire _guard91 = ev00__1_0;
wire _guard92 = ev00__1state >= 6'd1;
wire _guard93 = ev00__1state <= 6'd0;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = _guard91 | _guard94;
wire _guard96 = ev00__1_0;
wire _guard97 = ev00__1state >= 6'd1;
wire _guard98 = ev00__1state <= 6'd0;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = _guard96 | _guard99;
wire _guard101 = ev00__1_0;
wire _guard102 = ev00__1state >= 6'd1;
wire _guard103 = ev00__1state <= 6'd0;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = _guard101 | _guard104;
wire _guard106 = ev00__1_0;
wire _guard107 = ev00__1state >= 6'd1;
wire _guard108 = ev00__1state <= 6'd0;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = _guard106 | _guard109;
wire _guard111 = ev00__1_0;
wire _guard112 = ev00__1state >= 6'd1;
wire _guard113 = ev00__1state <= 6'd0;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = _guard111 | _guard114;
wire _guard116 = ev00__1_0;
wire _guard117 = ev00__1state >= 6'd1;
wire _guard118 = ev00__1state <= 6'd0;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = _guard116 | _guard119;
wire _guard121 = ev00__1_0;
wire _guard122 = ev00__1state >= 6'd1;
wire _guard123 = ev00__1state <= 6'd0;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = _guard121 | _guard124;
wire _guard126 = ev00__1_0;
wire _guard127 = ev00__1state >= 6'd1;
wire _guard128 = ev00__1state <= 6'd0;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = _guard126 | _guard129;
wire _guard131 = ev00__1_0;
wire _guard132 = ev00__1state >= 6'd1;
wire _guard133 = ev00__1state <= 6'd0;
wire _guard134 = _guard132 & _guard133;
wire _guard135 = _guard131 | _guard134;
wire _guard136 = ev00__1_0;
wire _guard137 = ev00__1state >= 6'd1;
wire _guard138 = ev00__1state <= 6'd0;
wire _guard139 = _guard137 & _guard138;
wire _guard140 = _guard136 | _guard139;
wire _guard141 = ev00__1_0;
wire _guard142 = ev00__1state >= 6'd1;
wire _guard143 = ev00__1state <= 6'd0;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = _guard141 | _guard144;
wire _guard146 = ev00__1_0;
wire _guard147 = ev00__1state >= 6'd1;
wire _guard148 = ev00__1state <= 6'd0;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = _guard146 | _guard149;
wire _guard151 = ev00__1_0;
wire _guard152 = ev00__1state >= 6'd1;
wire _guard153 = ev00__1state <= 6'd0;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = _guard151 | _guard154;
wire _guard156 = ev00__1_0;
wire _guard157 = ev00__1state >= 6'd1;
wire _guard158 = ev00__1state <= 6'd0;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = _guard156 | _guard159;
wire _guard161 = ev00__1_0;
wire _guard162 = ev00__1state >= 6'd1;
wire _guard163 = ev00__1state <= 6'd0;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = _guard161 | _guard164;
wire _guard166 = ev00__0_0;
wire _guard167 = ev00__0state >= 6'd1;
wire _guard168 = ev00__0state <= 6'd0;
wire _guard169 = _guard167 & _guard168;
wire _guard170 = _guard166 | _guard169;
wire _guard171 = ev00__0_0;
wire _guard172 = ev00__0state >= 6'd1;
wire _guard173 = ev00__0state <= 6'd0;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = _guard171 | _guard174;
wire _guard176 = ev00__0_0;
wire _guard177 = ev00__0state >= 6'd1;
wire _guard178 = ev00__0state <= 6'd0;
wire _guard179 = _guard177 & _guard178;
wire _guard180 = _guard176 | _guard179;
wire _guard181 = ev00__0_0;
wire _guard182 = ev00__0state >= 6'd1;
wire _guard183 = ev00__0state <= 6'd0;
wire _guard184 = _guard182 & _guard183;
wire _guard185 = _guard181 | _guard184;
wire _guard186 = ev00__0_0;
wire _guard187 = ev00__0state >= 6'd1;
wire _guard188 = ev00__0state <= 6'd0;
wire _guard189 = _guard187 & _guard188;
wire _guard190 = _guard186 | _guard189;
wire _guard191 = ev00__0_0;
wire _guard192 = ev00__0state >= 6'd1;
wire _guard193 = ev00__0state <= 6'd0;
wire _guard194 = _guard192 & _guard193;
wire _guard195 = _guard191 | _guard194;
wire _guard196 = ev00__0_0;
wire _guard197 = ev00__0state >= 6'd1;
wire _guard198 = ev00__0state <= 6'd0;
wire _guard199 = _guard197 & _guard198;
wire _guard200 = _guard196 | _guard199;
wire _guard201 = ev00__0_0;
wire _guard202 = ev00__0state >= 6'd1;
wire _guard203 = ev00__0state <= 6'd0;
wire _guard204 = _guard202 & _guard203;
wire _guard205 = _guard201 | _guard204;
wire _guard206 = ev00__0_0;
wire _guard207 = ev00__0state >= 6'd1;
wire _guard208 = ev00__0state <= 6'd0;
wire _guard209 = _guard207 & _guard208;
wire _guard210 = _guard206 | _guard209;
wire _guard211 = ev00__0_0;
wire _guard212 = ev00__0state >= 6'd1;
wire _guard213 = ev00__0state <= 6'd0;
wire _guard214 = _guard212 & _guard213;
wire _guard215 = _guard211 | _guard214;
wire _guard216 = ev00__0_0;
wire _guard217 = ev00__0state >= 6'd1;
wire _guard218 = ev00__0state <= 6'd0;
wire _guard219 = _guard217 & _guard218;
wire _guard220 = _guard216 | _guard219;
wire _guard221 = ev00__0_0;
wire _guard222 = ev00__0state >= 6'd1;
wire _guard223 = ev00__0state <= 6'd0;
wire _guard224 = _guard222 & _guard223;
wire _guard225 = _guard221 | _guard224;
wire _guard226 = ev00__0_0;
wire _guard227 = ev00__0state >= 6'd1;
wire _guard228 = ev00__0state <= 6'd0;
wire _guard229 = _guard227 & _guard228;
wire _guard230 = _guard226 | _guard229;
wire _guard231 = ev00__0_0;
wire _guard232 = ev00__0state >= 6'd1;
wire _guard233 = ev00__0state <= 6'd0;
wire _guard234 = _guard232 & _guard233;
wire _guard235 = _guard231 | _guard234;
wire _guard236 = ev00__0_0;
wire _guard237 = ev00__0state >= 6'd1;
wire _guard238 = ev00__0state <= 6'd0;
wire _guard239 = _guard237 & _guard238;
wire _guard240 = _guard236 | _guard239;
wire _guard241 = ev00__0_0;
wire _guard242 = ev00__0state >= 6'd1;
wire _guard243 = ev00__0state <= 6'd0;
wire _guard244 = _guard242 & _guard243;
wire _guard245 = _guard241 | _guard244;
wire _guard246 = ev00__0_0;
wire _guard247 = ev00__0state >= 6'd1;
wire _guard248 = ev00__0state <= 6'd0;
wire _guard249 = _guard247 & _guard248;
wire _guard250 = _guard246 | _guard249;
wire _guard251 = ev00__0_0;
wire _guard252 = ev00__0state >= 6'd1;
wire _guard253 = ev00__0state <= 6'd0;
wire _guard254 = _guard252 & _guard253;
wire _guard255 = _guard251 | _guard254;
wire _guard256 = ev00__0_0;
wire _guard257 = ev00__0state >= 6'd1;
wire _guard258 = ev00__0state <= 6'd0;
wire _guard259 = _guard257 & _guard258;
wire _guard260 = _guard256 | _guard259;
wire _guard261 = ev00__0_0;
wire _guard262 = ev00__0state >= 6'd1;
wire _guard263 = ev00__0state <= 6'd0;
wire _guard264 = _guard262 & _guard263;
wire _guard265 = _guard261 | _guard264;
wire _guard266 = ev00__0_0;
wire _guard267 = ev00__0state >= 6'd1;
wire _guard268 = ev00__0state <= 6'd0;
wire _guard269 = _guard267 & _guard268;
wire _guard270 = _guard266 | _guard269;
wire _guard271 = ev00__0_0;
wire _guard272 = ev00__0state >= 6'd1;
wire _guard273 = ev00__0state <= 6'd0;
wire _guard274 = _guard272 & _guard273;
wire _guard275 = _guard271 | _guard274;
wire _guard276 = ev00__0_0;
wire _guard277 = ev00__0state >= 6'd1;
wire _guard278 = ev00__0state <= 6'd0;
wire _guard279 = _guard277 & _guard278;
wire _guard280 = _guard276 | _guard279;
wire _guard281 = ev00__0_0;
wire _guard282 = ev00__0state >= 6'd1;
wire _guard283 = ev00__0state <= 6'd0;
wire _guard284 = _guard282 & _guard283;
wire _guard285 = _guard281 | _guard284;
wire _guard286 = ev00__0_0;
wire _guard287 = ev00__0state >= 6'd1;
wire _guard288 = ev00__0state <= 6'd0;
wire _guard289 = _guard287 & _guard288;
wire _guard290 = _guard286 | _guard289;
wire _guard291 = ev00__0_0;
wire _guard292 = ev00__0state >= 6'd1;
wire _guard293 = ev00__0state <= 6'd0;
wire _guard294 = _guard292 & _guard293;
wire _guard295 = _guard291 | _guard294;
wire _guard296 = ev00__0_0;
wire _guard297 = ev00__0state >= 6'd1;
wire _guard298 = ev00__0state <= 6'd0;
wire _guard299 = _guard297 & _guard298;
wire _guard300 = _guard296 | _guard299;
wire _guard301 = ev00__0_0;
wire _guard302 = ev00__0state >= 6'd1;
wire _guard303 = ev00__0state <= 6'd0;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = _guard301 | _guard304;
wire _guard306 = ev00__0_0;
wire _guard307 = ev00__0state >= 6'd1;
wire _guard308 = ev00__0state <= 6'd0;
wire _guard309 = _guard307 & _guard308;
wire _guard310 = _guard306 | _guard309;
wire _guard311 = ev00__0_0;
wire _guard312 = ev00__0state >= 6'd1;
wire _guard313 = ev00__0state <= 6'd0;
wire _guard314 = _guard312 & _guard313;
wire _guard315 = _guard311 | _guard314;
wire _guard316 = ev00__0_0;
wire _guard317 = ev00__0state >= 6'd1;
wire _guard318 = ev00__0state <= 6'd0;
wire _guard319 = _guard317 & _guard318;
wire _guard320 = _guard316 | _guard319;
wire _guard321 = ev00__0_0;
wire _guard322 = ev00__0state >= 6'd1;
wire _guard323 = ev00__0state <= 6'd0;
wire _guard324 = _guard322 & _guard323;
wire _guard325 = _guard321 | _guard324;
wire _guard326 = ev00__0_0;
wire _guard327 = ev00__0state >= 6'd1;
wire _guard328 = ev00__0state <= 6'd0;
wire _guard329 = _guard327 & _guard328;
wire _guard330 = _guard326 | _guard329;
assign p40 =
  _guard5 ? inst1_p39 :
  1024'd0;
assign inst1_p19 = inst0_p572;
assign inst1_p28 = inst0_p581;
assign inst1_p29 = inst0_p582;
assign inst1_p38 = inst0_p591;
assign inst1_p12 = inst0_p565;
assign inst1_p16 = inst0_p569;
assign inst1_p9 = inst0_p562;
assign inst1_p15 = inst0_p568;
assign inst1_p17 = inst0_p570;
assign inst1_p20 = inst0_p573;
assign inst1_p21 = inst0_p574;
assign inst1_p23 = inst0_p576;
assign inst1_clk = clk;
assign inst1_p11 = inst0_p564;
assign inst1_p25 = inst0_p578;
assign inst1_p36 = inst0_p589;
assign inst1_p8 = inst0_p561;
assign inst1_p10 = inst0_p563;
assign inst1_reset = reset;
assign inst1_p7 = inst0_p560;
assign inst1_p13 = inst0_p566;
assign inst1_p18 = inst0_p571;
assign inst1_p30 = inst0_p583;
assign inst1_p24 = inst0_p577;
assign inst1_p32 = inst0_p585;
assign inst1_p14 = inst0_p567;
assign inst1_p26 = inst0_p579;
assign inst1_p31 = inst0_p584;
assign inst1_p27 = inst0_p580;
assign inst1_p33 = inst0_p586;
assign inst1_p22 = inst0_p575;
assign inst1_p34 = inst0_p587;
assign inst1_p35 = inst0_p588;
assign inst1_p37 = inst0_p590;
assign inst0_ev0 = _guard170;
assign inst0_p533 = p13;
assign inst0_p559 = p39;
assign inst0_p534 = p14;
assign inst0_p556 = p36;
assign inst0_p540 = p20;
assign inst0_p551 = p31;
assign inst0_p537 = p17;
assign inst0_p542 = p22;
assign inst0_p545 = p25;
assign inst0_clk = clk;
assign inst0_p528 = p8;
assign inst0_p530 = p10;
assign inst0_p548 = p28;
assign inst0_p558 = p38;
assign inst0_p541 = p21;
assign inst0_p547 = p27;
assign inst0_p553 = p33;
assign inst0_p555 = p35;
assign inst0_p535 = p15;
assign inst0_p550 = p30;
assign inst0_reset = reset;
assign inst0_p536 = p16;
assign inst0_p544 = p24;
assign inst0_p546 = p26;
assign inst0_p538 = p18;
assign inst0_p554 = p34;
assign inst0_p557 = p37;
assign inst0_p543 = p23;
assign inst0_p552 = p32;
assign inst0_p529 = p9;
assign inst0_p549 = p29;
assign inst0_p539 = p19;
assign inst0_p532 = p12;
assign inst0_p531 = p11;
assign ev00_clk = clk;
assign ev00_go = ev0;
assign ev00_reset = reset;
// COMPONENT END: comp95
endmodule
module main(
  input logic [1023:0] in,
  output logic [1023:0] out,
  input logic go,
  input logic reset,
  input logic clk
);
// COMPONENT START: main
logic [5:0] go0__0state;
logic go0__0_0;
logic [5:0] go0__1state;
logic go0__1_0;
logic go0_clk;
logic go0_reset;
logic go0_go;
logic go0_done;
logic [1023:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [31:0] inst0_p38;
logic [31:0] inst0_p39;
logic [31:0] inst0_p40;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_p8;
logic [31:0] inst1_p9;
logic [31:0] inst1_p10;
logic [31:0] inst1_p11;
logic [31:0] inst1_p12;
logic [31:0] inst1_p13;
logic [31:0] inst1_p14;
logic [31:0] inst1_p15;
logic [31:0] inst1_p16;
logic [31:0] inst1_p17;
logic [31:0] inst1_p18;
logic [31:0] inst1_p19;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic [31:0] inst1_p30;
logic [31:0] inst1_p31;
logic [31:0] inst1_p32;
logic [31:0] inst1_p33;
logic [31:0] inst1_p34;
logic [31:0] inst1_p35;
logic [31:0] inst1_p36;
logic [31:0] inst1_p37;
logic [31:0] inst1_p38;
logic [31:0] inst1_p39;
logic [1023:0] inst1_p40;
logic inst1_ev0;
logic inst1_reset;
logic inst1_clk;
counter_chain_2_52 go0 (
    ._0_0(go0__0_0),
    ._0state(go0__0state),
    ._1_0(go0__1_0),
    ._1state(go0__1state),
    .clk(go0_clk),
    .done(go0_done),
    .go(go0_go),
    .reset(go0_reset)
);
comp32 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p39(inst0_p39),
    .p40(inst0_p40),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
comp95 inst1 (
    .clk(inst1_clk),
    .ev0(inst1_ev0),
    .p10(inst1_p10),
    .p11(inst1_p11),
    .p12(inst1_p12),
    .p13(inst1_p13),
    .p14(inst1_p14),
    .p15(inst1_p15),
    .p16(inst1_p16),
    .p17(inst1_p17),
    .p18(inst1_p18),
    .p19(inst1_p19),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .p30(inst1_p30),
    .p31(inst1_p31),
    .p32(inst1_p32),
    .p33(inst1_p33),
    .p34(inst1_p34),
    .p35(inst1_p35),
    .p36(inst1_p36),
    .p37(inst1_p37),
    .p38(inst1_p38),
    .p39(inst1_p39),
    .p40(inst1_p40),
    .p8(inst1_p8),
    .p9(inst1_p9),
    .reset(inst1_reset)
);
wire _guard0 = 1;
wire _guard1 = go0__1_0;
wire _guard2 = go0__1state >= 6'd1;
wire _guard3 = go0__1state <= 6'd0;
wire _guard4 = _guard2 & _guard3;
wire _guard5 = _guard1 | _guard4;
wire _guard6 = go0__0_0;
wire _guard7 = go0__0state >= 6'd1;
wire _guard8 = go0__0state <= 6'd0;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = _guard6 | _guard9;
wire _guard11 = go0__0_0;
wire _guard12 = go0__0state >= 6'd1;
wire _guard13 = go0__0state <= 6'd0;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = _guard11 | _guard14;
wire _guard16 = go0__0_0;
wire _guard17 = go0__0state >= 6'd1;
wire _guard18 = go0__0state <= 6'd0;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = _guard16 | _guard19;
wire _guard21 = go0__0_0;
wire _guard22 = go0__0state >= 6'd1;
wire _guard23 = go0__0state <= 6'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard21 | _guard24;
wire _guard26 = go0__0_0;
wire _guard27 = go0__0state >= 6'd1;
wire _guard28 = go0__0state <= 6'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard26 | _guard29;
wire _guard31 = go0__0_0;
wire _guard32 = go0__0state >= 6'd1;
wire _guard33 = go0__0state <= 6'd0;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = _guard31 | _guard34;
wire _guard36 = go0__0_0;
wire _guard37 = go0__0state >= 6'd1;
wire _guard38 = go0__0state <= 6'd0;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = _guard36 | _guard39;
wire _guard41 = go0__0_0;
wire _guard42 = go0__0state >= 6'd1;
wire _guard43 = go0__0state <= 6'd0;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = _guard41 | _guard44;
wire _guard46 = go0__0_0;
wire _guard47 = go0__0state >= 6'd1;
wire _guard48 = go0__0state <= 6'd0;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = _guard46 | _guard49;
wire _guard51 = go0__0_0;
wire _guard52 = go0__0state >= 6'd1;
wire _guard53 = go0__0state <= 6'd0;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = _guard51 | _guard54;
wire _guard56 = go0__0_0;
wire _guard57 = go0__0state >= 6'd1;
wire _guard58 = go0__0state <= 6'd0;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = _guard56 | _guard59;
wire _guard61 = go0__0_0;
wire _guard62 = go0__0state >= 6'd1;
wire _guard63 = go0__0state <= 6'd0;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = _guard61 | _guard64;
wire _guard66 = go0__0_0;
wire _guard67 = go0__0state >= 6'd1;
wire _guard68 = go0__0state <= 6'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = _guard66 | _guard69;
wire _guard71 = go0__0_0;
wire _guard72 = go0__0state >= 6'd1;
wire _guard73 = go0__0state <= 6'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard71 | _guard74;
wire _guard76 = go0__0_0;
wire _guard77 = go0__0state >= 6'd1;
wire _guard78 = go0__0state <= 6'd0;
wire _guard79 = _guard77 & _guard78;
wire _guard80 = _guard76 | _guard79;
wire _guard81 = go0__0_0;
wire _guard82 = go0__0state >= 6'd1;
wire _guard83 = go0__0state <= 6'd0;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = _guard81 | _guard84;
wire _guard86 = go0__0_0;
wire _guard87 = go0__0state >= 6'd1;
wire _guard88 = go0__0state <= 6'd0;
wire _guard89 = _guard87 & _guard88;
wire _guard90 = _guard86 | _guard89;
wire _guard91 = go0__0_0;
wire _guard92 = go0__0state >= 6'd1;
wire _guard93 = go0__0state <= 6'd0;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = _guard91 | _guard94;
wire _guard96 = go0__0_0;
wire _guard97 = go0__0state >= 6'd1;
wire _guard98 = go0__0state <= 6'd0;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = _guard96 | _guard99;
wire _guard101 = go0__0_0;
wire _guard102 = go0__0state >= 6'd1;
wire _guard103 = go0__0state <= 6'd0;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = _guard101 | _guard104;
wire _guard106 = go0__0_0;
wire _guard107 = go0__0state >= 6'd1;
wire _guard108 = go0__0state <= 6'd0;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = _guard106 | _guard109;
wire _guard111 = go0__0_0;
wire _guard112 = go0__0state >= 6'd1;
wire _guard113 = go0__0state <= 6'd0;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = _guard111 | _guard114;
wire _guard116 = go0__0_0;
wire _guard117 = go0__0state >= 6'd1;
wire _guard118 = go0__0state <= 6'd0;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = _guard116 | _guard119;
wire _guard121 = go0__0_0;
wire _guard122 = go0__0state >= 6'd1;
wire _guard123 = go0__0state <= 6'd0;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = _guard121 | _guard124;
wire _guard126 = go0__0_0;
wire _guard127 = go0__0state >= 6'd1;
wire _guard128 = go0__0state <= 6'd0;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = _guard126 | _guard129;
wire _guard131 = go0__0_0;
wire _guard132 = go0__0state >= 6'd1;
wire _guard133 = go0__0state <= 6'd0;
wire _guard134 = _guard132 & _guard133;
wire _guard135 = _guard131 | _guard134;
wire _guard136 = go0__0_0;
wire _guard137 = go0__0state >= 6'd1;
wire _guard138 = go0__0state <= 6'd0;
wire _guard139 = _guard137 & _guard138;
wire _guard140 = _guard136 | _guard139;
wire _guard141 = go0__0_0;
wire _guard142 = go0__0state >= 6'd1;
wire _guard143 = go0__0state <= 6'd0;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = _guard141 | _guard144;
wire _guard146 = go0__0_0;
wire _guard147 = go0__0state >= 6'd1;
wire _guard148 = go0__0state <= 6'd0;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = _guard146 | _guard149;
wire _guard151 = go0__0_0;
wire _guard152 = go0__0state >= 6'd1;
wire _guard153 = go0__0state <= 6'd0;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = _guard151 | _guard154;
wire _guard156 = go0__0_0;
wire _guard157 = go0__0state >= 6'd1;
wire _guard158 = go0__0state <= 6'd0;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = _guard156 | _guard159;
wire _guard161 = go0__0_0;
wire _guard162 = go0__0state >= 6'd1;
wire _guard163 = go0__0state <= 6'd0;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = _guard161 | _guard164;
wire _guard166 = go0__0_0;
wire _guard167 = go0__0state >= 6'd1;
wire _guard168 = go0__0state <= 6'd0;
wire _guard169 = _guard167 & _guard168;
wire _guard170 = _guard166 | _guard169;
wire _guard171 = go0__0_0;
wire _guard172 = go0__0state >= 6'd1;
wire _guard173 = go0__0state <= 6'd0;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = _guard171 | _guard174;
assign out =
  _guard5 ? inst1_p40 :
  1024'd0;
assign go0_clk = clk;
assign go0_go = go;
assign go0_reset = reset;
assign inst1_p19 = inst0_p20;
assign inst1_p28 = inst0_p29;
assign inst1_p29 = inst0_p30;
assign inst1_p38 = inst0_p39;
assign inst1_p12 = inst0_p13;
assign inst1_p16 = inst0_p17;
assign inst1_ev0 = _guard40;
assign inst1_p9 = inst0_p10;
assign inst1_p15 = inst0_p16;
assign inst1_p17 = inst0_p18;
assign inst1_p20 = inst0_p21;
assign inst1_p21 = inst0_p22;
assign inst1_p23 = inst0_p24;
assign inst1_clk = clk;
assign inst1_p11 = inst0_p12;
assign inst1_p25 = inst0_p26;
assign inst1_p36 = inst0_p37;
assign inst1_p39 = inst0_p40;
assign inst1_p8 = inst0_p9;
assign inst1_p10 = inst0_p11;
assign inst1_reset = reset;
assign inst1_p13 = inst0_p14;
assign inst1_p18 = inst0_p19;
assign inst1_p30 = inst0_p31;
assign inst1_p24 = inst0_p25;
assign inst1_p32 = inst0_p33;
assign inst1_p14 = inst0_p15;
assign inst1_p26 = inst0_p27;
assign inst1_p31 = inst0_p32;
assign inst1_p27 = inst0_p28;
assign inst1_p33 = inst0_p34;
assign inst1_p22 = inst0_p23;
assign inst1_p34 = inst0_p35;
assign inst1_p35 = inst0_p36;
assign inst1_p37 = inst0_p38;
assign inst0_clk = clk;
assign inst0_p8 = in;
assign inst0_reset = reset;
// COMPONENT END: main
endmodule
module counter_52(
  input logic clk,
  input logic reset,
  output logic [5:0] state,
  output logic _0,
  input logic go,
  output logic done
);
// COMPONENT START: counter_52
logic [5:0] add_left;
logic [5:0] add_right;
logic [5:0] add_out;
logic [5:0] state0_in;
logic state0_write_en;
logic state0_clk;
logic state0_reset;
logic [5:0] state0_out;
logic state0_done;
logic done0_in;
logic done0_write_en;
logic done0_clk;
logic done0_reset;
logic done0_out;
logic done0_done;
std_add # (
    .WIDTH(6)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
std_reg # (
    .WIDTH(6)
) state0 (
    .clk(state0_clk),
    .done(state0_done),
    .in(state0_in),
    .out(state0_out),
    .reset(state0_reset),
    .write_en(state0_write_en)
);
std_reg # (
    .WIDTH(1)
) done0 (
    .clk(done0_clk),
    .done(done0_done),
    .in(done0_in),
    .out(done0_out),
    .reset(done0_reset),
    .write_en(done0_write_en)
);
wire _guard0 = 1;
wire _guard1 = go;
wire _guard2 = state0_out == 6'd0;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = state0_out == 6'd51;
wire _guard5 = state0_out != 6'd51;
wire _guard6 = state0_out == 6'd51;
wire _guard7 = go;
wire _guard8 = state0_out != 6'd0;
wire _guard9 = _guard7 | _guard8;
wire _guard10 = state0_out != 6'd51;
wire _guard11 = _guard9 & _guard10;
wire _guard12 = _guard6 | _guard11;
wire _guard13 = state0_out == 6'd51;
wire _guard14 = go;
wire _guard15 = state0_out != 6'd0;
wire _guard16 = _guard14 | _guard15;
wire _guard17 = state0_out != 6'd51;
wire _guard18 = _guard16 & _guard17;
assign done = done0_out;
assign _0 = _guard3;
assign state = state0_out;
assign add_left = state0_out;
assign add_right = 6'd1;
assign done0_write_en = 1'd1;
assign done0_clk = clk;
assign done0_reset = reset;
assign done0_in =
  _guard4 ? 1'd1 :
  _guard5 ? 1'd0 :
  'x;
assign state0_write_en = _guard12;
assign state0_clk = clk;
assign state0_reset = reset;
assign state0_in =
  _guard13 ? 6'd0 :
  _guard18 ? add_out :
  'x;
// COMPONENT END: counter_52
endmodule
module fsm_5(
  output logic _0,
  output logic _1,
  output logic _2,
  output logic _3,
  output logic _4,
  input logic clk,
  input logic reset,
  input logic go,
  output logic done
);
// COMPONENT START: fsm_5
logic r_in;
logic r_write_en;
logic r_clk;
logic r_reset;
logic r_out;
logic r_done;
logic r0_in;
logic r0_write_en;
logic r0_clk;
logic r0_reset;
logic r0_out;
logic r0_done;
logic r1_in;
logic r1_write_en;
logic r1_clk;
logic r1_reset;
logic r1_out;
logic r1_done;
logic r2_in;
logic r2_write_en;
logic r2_clk;
logic r2_reset;
logic r2_out;
logic r2_done;
logic r3_in;
logic r3_write_en;
logic r3_clk;
logic r3_reset;
logic r3_out;
logic r3_done;
std_reg # (
    .WIDTH(1)
) r (
    .clk(r_clk),
    .done(r_done),
    .in(r_in),
    .out(r_out),
    .reset(r_reset),
    .write_en(r_write_en)
);
std_reg # (
    .WIDTH(1)
) r0 (
    .clk(r0_clk),
    .done(r0_done),
    .in(r0_in),
    .out(r0_out),
    .reset(r0_reset),
    .write_en(r0_write_en)
);
std_reg # (
    .WIDTH(1)
) r1 (
    .clk(r1_clk),
    .done(r1_done),
    .in(r1_in),
    .out(r1_out),
    .reset(r1_reset),
    .write_en(r1_write_en)
);
std_reg # (
    .WIDTH(1)
) r2 (
    .clk(r2_clk),
    .done(r2_done),
    .in(r2_in),
    .out(r2_out),
    .reset(r2_reset),
    .write_en(r2_write_en)
);
std_reg # (
    .WIDTH(1)
) r3 (
    .clk(r3_clk),
    .done(r3_done),
    .in(r3_in),
    .out(r3_out),
    .reset(r3_reset),
    .write_en(r3_write_en)
);
wire _guard0 = 1;
assign done = r3_out;
assign _2 = r0_out;
assign _1 = r_out;
assign _0 = go;
assign _3 = r1_out;
assign _4 = r2_out;
assign r_write_en = 1'd1;
assign r_clk = clk;
assign r_reset = reset;
assign r_in = go;
assign r0_write_en = 1'd1;
assign r0_clk = clk;
assign r0_reset = reset;
assign r0_in = r_out;
assign r1_write_en = 1'd1;
assign r1_clk = clk;
assign r1_reset = reset;
assign r1_in = r0_out;
assign r2_write_en = 1'd1;
assign r2_clk = clk;
assign r2_reset = reset;
assign r2_in = r1_out;
assign r3_write_en = 1'd1;
assign r3_clk = clk;
assign r3_reset = reset;
assign r3_in = r2_out;
// COMPONENT END: fsm_5
endmodule
module counter_chain_2_52(
  output logic [5:0] _0state,
  output logic _0_0,
  output logic [5:0] _1state,
  output logic _1_0,
  input logic clk,
  input logic reset,
  input logic go,
  output logic done
);
// COMPONENT START: counter_chain_2_52
logic c0_clk;
logic c0_reset;
logic [5:0] c0_state;
logic c0__0;
logic c0_go;
logic c0_done;
logic c1_clk;
logic c1_reset;
logic [5:0] c1_state;
logic c1__0;
logic c1_go;
logic c1_done;
counter_52 c0 (
    ._0(c0__0),
    .clk(c0_clk),
    .done(c0_done),
    .go(c0_go),
    .reset(c0_reset),
    .state(c0_state)
);
counter_52 c1 (
    ._0(c1__0),
    .clk(c1_clk),
    .done(c1_done),
    .go(c1_go),
    .reset(c1_reset),
    .state(c1_state)
);
wire _guard0 = 1;
assign done = c1_done;
assign _0state = c0_state;
assign _1state = c1_state;
assign _0_0 = c0__0;
assign _1_0 = c1__0;
assign c1_clk = clk;
assign c1_go = c0_done;
assign c1_reset = reset;
assign c0_clk = clk;
assign c0_go = go;
assign c0_reset = reset;
// COMPONENT END: counter_chain_2_52
endmodule
