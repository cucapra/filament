module Neg #(
  parameter WIDTH = 32
) (
  input wire logic signed [WIDTH-1:0] in,
  output wire logic signed [WIDTH-1:0] out
);
  assign out = -in;
endmodule
`default_nettype none

module Register #(
    parameter WIDTH = 32
) (
  input wire clk,
  input wire reset,
  input wire logic write_en,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] out
);
  always_ff @(posedge clk) begin
    if (reset)
      out <= 0;
    else if (write_en)
      out <= in;
    else
      out <= out;
  end
endmodule

// Same as a register but does not have a write enable signal.
module Delay #(
    parameter WIDTH = 32
) (
  input wire clk,
  input wire reset,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] out
);

  Register #(WIDTH) r (
    .clk(clk),
    .reset(reset),
    .write_en(1'b1),
    .in(in),
    .out(out)
  );
endmodule

// Register that passes its input value through.
module PassThroughRegister #(
  parameter WIDTH = 32
) (
  input wire clk,
  input wire reset,
  input wire logic write_en,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] out
);
  // held register value
  logic [WIDTH-1:0] t_out;
  Register #(WIDTH) r (
    .clk(clk),
    .reset(reset),
    .write_en(write_en),
    .in(in),
    .out(t_out)
  );
  
  assign out = write_en ? in : t_out;
endmodule

// Similar to a register but provides access to its previous value only.
// Resetting behavior controlled using the SAFE parameter.
module Prev #(
    parameter WIDTH = 32,
    // If 0, reset to 'x, otherwise reset to 0
    parameter SAFE = 0
) (
  input wire clk,
  input wire reset,
  input wire logic write_en,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] prev
);
  always_ff @(posedge clk) begin
    if (reset)
      if (SAFE == 0)
        prev <= 'x;
      else
        prev <= '0;
    else if (write_en)
      prev <= in;
    else
      prev <= prev;
  end
endmodule

module ContPrev #(
    parameter WIDTH = 32,
    parameter SAFE = 0
) (
  input wire clk,
  input wire reset,
  input wire logic [WIDTH-1:0] in,
  output logic [WIDTH-1:0] prev
);

Prev #(WIDTH, SAFE) r (
  .clk(clk),
  .reset(reset),
  .write_en(1'b1),
  .in(in),
  .prev(prev)
);
endmodule


`default_nettype wire
module Butterfly_Exp8_Mant23(
  input wire clk,
  input wire [31:0] in0_r,
  input wire [31:0] in0_i,
  input wire [31:0] in1_r,
  input wire [31:0] in1_i,
  input wire [31:0] twd_r,
  input wire [31:0] twd_i,
  output wire [127:0] out
);
  // lint_off MULTIPLY
  function automatic [47:0] umul48b_24b_x_24b (input reg [23:0] lhs, input reg [23:0] rhs);
    begin
      umul48b_24b_x_24b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY

  // ===== Pipe stage 0:
  wire [2:0] p0_literal_8123_comb;
  wire [2:0] p0_literal_8129_comb;
  wire [2:0] p0_literal_8134_comb;
  wire [2:0] p0_literal_8140_comb;
  assign p0_literal_8123_comb = 3'h0;
  assign p0_literal_8129_comb = 3'h0;
  assign p0_literal_8134_comb = 3'h0;
  assign p0_literal_8140_comb = 3'h0;

  // Registers for pipe stage 0:
  reg [31:0] p0_in0_r;
  reg [31:0] p0_in0_i;
  reg [31:0] p0_in1_r;
  reg [31:0] p0_in1_i;
  reg [31:0] p0_twd_r;
  reg [31:0] p0_twd_i;
  reg [2:0] p7_literal_8123;
  reg [2:0] p7_literal_8129;
  reg [2:0] p7_literal_8134;
  reg [2:0] p7_literal_8140;
  always_ff @ (posedge clk) begin
    p0_in0_r <= in0_r;
    p0_in0_i <= in0_i;
    p0_in1_r <= in1_r;
    p0_in1_i <= in1_i;
    p0_twd_r <= twd_r;
    p0_twd_i <= twd_i;
    p7_literal_8123 <= p0_literal_8123_comb;
    p7_literal_8129 <= p0_literal_8129_comb;
    p7_literal_8134 <= p0_literal_8134_comb;
    p7_literal_8140 <= p0_literal_8140_comb;
  end

  // ===== Pipe stage 1:
  wire [22:0] p1_in1_r_fraction__10_comb;
  wire [7:0] p1_in1_r_bexp__9_comb;
  wire [22:0] p1_twd_r_fraction__10_comb;
  wire [7:0] p1_twd_r_bexp__9_comb;
  wire [22:0] p1_in1_i_fraction__10_comb;
  wire [7:0] p1_in1_i_bexp__9_comb;
  wire [22:0] p1_twd_i_fraction__10_comb;
  wire [7:0] p1_twd_i_bexp__9_comb;
  wire [7:0] p1_high_exp__3_comb;
  wire [7:0] p1_high_exp__4_comb;
  wire [7:0] p1_high_exp__6_comb;
  wire [7:0] p1_high_exp__1_comb;
  wire [23:0] p1_in1_r_fraction__11_comb;
  wire [23:0] p1_twd_r_fraction__11_comb;
  wire [23:0] p1_in1_i_fraction__11_comb;
  wire [23:0] p1_twd_i_fraction__11_comb;
  wire [8:0] p1_concat_7295_comb;
  wire [8:0] p1_concat_7296_comb;
  wire [8:0] p1_concat_7301_comb;
  wire [8:0] p1_concat_7302_comb;
  wire p1_eq_7323_comb;
  wire p1_eq_7325_comb;
  wire p1_eq_7327_comb;
  wire p1_eq_7329_comb;
  wire p1_in1_i_sign__2_comb;
  wire p1_twd_i_sign__2_comb;
  wire p1_in1_r_sign__2_comb;
  wire p1_twd_r_sign__2_comb;
  wire [23:0] p1_in1_r_fraction__12_comb;
  wire [23:0] p1_twd_r_fraction__12_comb;
  wire [23:0] p1_in1_i_fraction__12_comb;
  wire [23:0] p1_twd_i_fraction__12_comb;
  wire [8:0] p1_add_7307_comb;
  wire p1_eq_7308_comb;
  wire p1_eq_7309_comb;
  wire [8:0] p1_add_7310_comb;
  wire p1_eq_7311_comb;
  wire p1_eq_7312_comb;
  wire [8:0] p1_add_7313_comb;
  wire [8:0] p1_add_7314_comb;
  wire p1_and_7333_comb;
  wire p1_and_7334_comb;
  wire p1_and_7337_comb;
  wire p1_and_7338_comb;
  wire p1_and_7343_comb;
  wire p1_and_7344_comb;
  wire p1_and_7345_comb;
  wire p1_and_7346_comb;
  wire p1_result_sign__2_comb;
  wire p1_result_sign__1_comb;
  wire p1_result_sign__6_comb;
  wire p1_result_sign__4_comb;
  wire [22:0] p1_in0_r_fraction__6_comb;
  wire [7:0] p1_in0_r_bexp__6_comb;
  wire [22:0] p1_in0_i_fraction__6_comb;
  wire [7:0] p1_in0_i_bexp__6_comb;
  wire p1_in0_r_sign__2_comb;
  wire p1_in0_i_sign__2_comb;
  assign p1_in1_r_fraction__10_comb = p0_in1_r[22:0];
  assign p1_in1_r_bexp__9_comb = p0_in1_r[30:23];
  assign p1_twd_r_fraction__10_comb = p0_twd_r[22:0];
  assign p1_twd_r_bexp__9_comb = p0_twd_r[30:23];
  assign p1_in1_i_fraction__10_comb = p0_in1_i[22:0];
  assign p1_in1_i_bexp__9_comb = p0_in1_i[30:23];
  assign p1_twd_i_fraction__10_comb = p0_twd_i[22:0];
  assign p1_twd_i_bexp__9_comb = p0_twd_i[30:23];
  assign p1_high_exp__3_comb = 8'hff;
  assign p1_high_exp__4_comb = 8'hff;
  assign p1_high_exp__6_comb = 8'hff;
  assign p1_high_exp__1_comb = 8'hff;
  assign p1_in1_r_fraction__11_comb = {1'h0, p1_in1_r_fraction__10_comb} | 24'h80_0000;
  assign p1_twd_r_fraction__11_comb = {1'h0, p1_twd_r_fraction__10_comb} | 24'h80_0000;
  assign p1_in1_i_fraction__11_comb = {1'h0, p1_in1_i_fraction__10_comb} | 24'h80_0000;
  assign p1_twd_i_fraction__11_comb = {1'h0, p1_twd_i_fraction__10_comb} | 24'h80_0000;
  assign p1_concat_7295_comb = {1'h0, p1_in1_r_bexp__9_comb};
  assign p1_concat_7296_comb = {1'h0, p1_twd_r_bexp__9_comb};
  assign p1_concat_7301_comb = {1'h0, p1_in1_i_bexp__9_comb};
  assign p1_concat_7302_comb = {1'h0, p1_twd_i_bexp__9_comb};
  assign p1_eq_7323_comb = p1_in1_r_bexp__9_comb == p1_high_exp__3_comb;
  assign p1_eq_7325_comb = p1_twd_r_bexp__9_comb == p1_high_exp__4_comb;
  assign p1_eq_7327_comb = p1_in1_i_bexp__9_comb == p1_high_exp__6_comb;
  assign p1_eq_7329_comb = p1_twd_i_bexp__9_comb == p1_high_exp__1_comb;
  assign p1_in1_i_sign__2_comb = p0_in1_i[31:31];
  assign p1_twd_i_sign__2_comb = p0_twd_i[31:31];
  assign p1_in1_r_sign__2_comb = p0_in1_r[31:31];
  assign p1_twd_r_sign__2_comb = p0_twd_r[31:31];
  assign p1_in1_r_fraction__12_comb = p1_in1_r_fraction__11_comb & {24{p1_in1_r_bexp__9_comb != 8'h00}};
  assign p1_twd_r_fraction__12_comb = p1_twd_r_fraction__11_comb & {24{p1_twd_r_bexp__9_comb != 8'h00}};
  assign p1_in1_i_fraction__12_comb = p1_in1_i_fraction__11_comb & {24{p1_in1_i_bexp__9_comb != 8'h00}};
  assign p1_twd_i_fraction__12_comb = p1_twd_i_fraction__11_comb & {24{p1_twd_i_bexp__9_comb != 8'h00}};
  assign p1_add_7307_comb = p1_concat_7295_comb + p1_concat_7296_comb;
  assign p1_eq_7308_comb = p1_in1_r_bexp__9_comb == 8'h00;
  assign p1_eq_7309_comb = p1_twd_r_bexp__9_comb == 8'h00;
  assign p1_add_7310_comb = p1_concat_7301_comb + p1_concat_7302_comb;
  assign p1_eq_7311_comb = p1_in1_i_bexp__9_comb == 8'h00;
  assign p1_eq_7312_comb = p1_twd_i_bexp__9_comb == 8'h00;
  assign p1_add_7313_comb = p1_concat_7295_comb + p1_concat_7302_comb;
  assign p1_add_7314_comb = p1_concat_7301_comb + p1_concat_7296_comb;
  assign p1_and_7333_comb = p1_eq_7323_comb & p1_in1_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_7334_comb = p1_eq_7325_comb & p1_twd_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_7337_comb = p1_eq_7327_comb & p1_in1_i_fraction__10_comb == 23'h00_0000;
  assign p1_and_7338_comb = p1_eq_7329_comb & p1_twd_i_fraction__10_comb == 23'h00_0000;
  assign p1_and_7343_comb = p1_eq_7323_comb & p1_in1_r_fraction__10_comb != 23'h00_0000;
  assign p1_and_7344_comb = p1_eq_7325_comb & p1_twd_r_fraction__10_comb != 23'h00_0000;
  assign p1_and_7345_comb = p1_eq_7327_comb & p1_in1_i_fraction__10_comb != 23'h00_0000;
  assign p1_and_7346_comb = p1_eq_7329_comb & p1_twd_i_fraction__10_comb != 23'h00_0000;
  assign p1_result_sign__2_comb = p1_in1_i_sign__2_comb ^ p1_twd_i_sign__2_comb;
  assign p1_result_sign__1_comb = p1_in1_r_sign__2_comb ^ p1_twd_r_sign__2_comb;
  assign p1_result_sign__6_comb = p1_in1_i_sign__2_comb ^ p1_twd_r_sign__2_comb;
  assign p1_result_sign__4_comb = p1_in1_r_sign__2_comb ^ p1_twd_i_sign__2_comb;
  assign p1_in0_r_fraction__6_comb = p0_in0_r[22:0];
  assign p1_in0_r_bexp__6_comb = p0_in0_r[30:23];
  assign p1_in0_i_fraction__6_comb = p0_in0_i[22:0];
  assign p1_in0_i_bexp__6_comb = p0_in0_i[30:23];
  assign p1_in0_r_sign__2_comb = p0_in0_r[31:31];
  assign p1_in0_i_sign__2_comb = p0_in0_i[31:31];

  // Registers for pipe stage 1:
  reg [23:0] p1_in1_r_fraction__12;
  reg [23:0] p1_twd_r_fraction__12;
  reg [23:0] p1_in1_i_fraction__12;
  reg [23:0] p1_twd_i_fraction__12;
  reg [8:0] p1_add_7307;
  reg p1_eq_7308;
  reg p1_eq_7309;
  reg [8:0] p1_add_7310;
  reg p1_eq_7311;
  reg p1_eq_7312;
  reg [8:0] p1_add_7313;
  reg [8:0] p1_add_7314;
  reg p1_and_7333;
  reg p1_and_7334;
  reg p1_and_7337;
  reg p1_and_7338;
  reg p1_and_7343;
  reg p1_and_7344;
  reg p1_and_7345;
  reg p1_and_7346;
  reg p1_result_sign__2;
  reg p1_result_sign__1;
  reg p1_result_sign__6;
  reg p1_result_sign__4;
  reg [22:0] p1_in0_r_fraction__6;
  reg [7:0] p1_in0_r_bexp__6;
  reg [22:0] p1_in0_i_fraction__6;
  reg [7:0] p1_in0_i_bexp__6;
  reg p1_in0_r_sign__2;
  reg p1_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p1_in1_r_fraction__12 <= p1_in1_r_fraction__12_comb;
    p1_twd_r_fraction__12 <= p1_twd_r_fraction__12_comb;
    p1_in1_i_fraction__12 <= p1_in1_i_fraction__12_comb;
    p1_twd_i_fraction__12 <= p1_twd_i_fraction__12_comb;
    p1_add_7307 <= p1_add_7307_comb;
    p1_eq_7308 <= p1_eq_7308_comb;
    p1_eq_7309 <= p1_eq_7309_comb;
    p1_add_7310 <= p1_add_7310_comb;
    p1_eq_7311 <= p1_eq_7311_comb;
    p1_eq_7312 <= p1_eq_7312_comb;
    p1_add_7313 <= p1_add_7313_comb;
    p1_add_7314 <= p1_add_7314_comb;
    p1_and_7333 <= p1_and_7333_comb;
    p1_and_7334 <= p1_and_7334_comb;
    p1_and_7337 <= p1_and_7337_comb;
    p1_and_7338 <= p1_and_7338_comb;
    p1_and_7343 <= p1_and_7343_comb;
    p1_and_7344 <= p1_and_7344_comb;
    p1_and_7345 <= p1_and_7345_comb;
    p1_and_7346 <= p1_and_7346_comb;
    p1_result_sign__2 <= p1_result_sign__2_comb;
    p1_result_sign__1 <= p1_result_sign__1_comb;
    p1_result_sign__6 <= p1_result_sign__6_comb;
    p1_result_sign__4 <= p1_result_sign__4_comb;
    p1_in0_r_fraction__6 <= p1_in0_r_fraction__6_comb;
    p1_in0_r_bexp__6 <= p1_in0_r_bexp__6_comb;
    p1_in0_i_fraction__6 <= p1_in0_i_fraction__6_comb;
    p1_in0_i_bexp__6 <= p1_in0_i_bexp__6_comb;
    p1_in0_r_sign__2 <= p1_in0_r_sign__2_comb;
    p1_in0_i_sign__2 <= p1_in0_i_sign__2_comb;
  end

  // ===== Pipe stage 2:
  wire p2_has_0_arg__1_comb;
  wire p2_has_inf_arg__1_comb;
  wire p2_has_0_arg__2_comb;
  wire p2_has_inf_arg__2_comb;
  wire p2_has_0_arg__4_comb;
  wire p2_has_inf_arg__4_comb;
  wire p2_has_0_arg__3_comb;
  wire p2_has_inf_arg__3_comb;
  wire [47:0] p2_fraction__1_comb;
  wire [47:0] p2_fraction__8_comb;
  wire [47:0] p2_fraction__16_comb;
  wire [47:0] p2_fraction__24_comb;
  wire [9:0] p2_exp__1_comb;
  wire [9:0] p2_exp__4_comb;
  wire [9:0] p2_exp__8_comb;
  wire [9:0] p2_exp__12_comb;
  wire p2_is_result_nan__1_comb;
  wire p2_is_result_nan__2_comb;
  wire p2_is_result_nan__4_comb;
  wire p2_is_result_nan__3_comb;
  wire [47:0] p2_fraction__2_comb;
  wire [47:0] p2_sticky__1_comb;
  wire [47:0] p2_fraction__9_comb;
  wire [47:0] p2_sticky__2_comb;
  wire [47:0] p2_fraction__17_comb;
  wire [47:0] p2_sticky__4_comb;
  wire [47:0] p2_fraction__25_comb;
  wire [47:0] p2_sticky__6_comb;
  wire [9:0] p2_exp__2_comb;
  wire [9:0] p2_exp__5_comb;
  wire [9:0] p2_exp__9_comb;
  wire [9:0] p2_exp__13_comb;
  wire [47:0] p2_fraction__3_comb;
  wire [47:0] p2_fraction__10_comb;
  wire [47:0] p2_fraction__18_comb;
  wire [47:0] p2_fraction__26_comb;
  wire [9:0] p2_exp__3_comb;
  wire [9:0] p2_exp__6_comb;
  wire [9:0] p2_exp__10_comb;
  wire [9:0] p2_exp__14_comb;
  wire p2_nor_7497_comb;
  wire p2_nor_7499_comb;
  wire p2_nor_7501_comb;
  wire p2_nor_7503_comb;
  wire p2_result_sign__3_comb;
  wire p2_result_sign__5_comb;
  wire p2_result_sign__8_comb;
  wire p2_result_sign__7_comb;
  assign p2_has_0_arg__1_comb = p1_eq_7311 | p1_eq_7312;
  assign p2_has_inf_arg__1_comb = p1_and_7337 | p1_and_7338;
  assign p2_has_0_arg__2_comb = p1_eq_7308 | p1_eq_7309;
  assign p2_has_inf_arg__2_comb = p1_and_7333 | p1_and_7334;
  assign p2_has_0_arg__4_comb = p1_eq_7311 | p1_eq_7309;
  assign p2_has_inf_arg__4_comb = p1_and_7337 | p1_and_7334;
  assign p2_has_0_arg__3_comb = p1_eq_7308 | p1_eq_7312;
  assign p2_has_inf_arg__3_comb = p1_and_7333 | p1_and_7338;
  assign p2_fraction__1_comb = umul48b_24b_x_24b(p1_in1_r_fraction__12, p1_twd_r_fraction__12);
  assign p2_fraction__8_comb = umul48b_24b_x_24b(p1_in1_i_fraction__12, p1_twd_i_fraction__12);
  assign p2_fraction__16_comb = umul48b_24b_x_24b(p1_in1_r_fraction__12, p1_twd_i_fraction__12);
  assign p2_fraction__24_comb = umul48b_24b_x_24b(p1_in1_i_fraction__12, p1_twd_r_fraction__12);
  assign p2_exp__1_comb = {1'h0, p1_add_7307} + 10'h381;
  assign p2_exp__4_comb = {1'h0, p1_add_7310} + 10'h381;
  assign p2_exp__8_comb = {1'h0, p1_add_7313} + 10'h381;
  assign p2_exp__12_comb = {1'h0, p1_add_7314} + 10'h381;
  assign p2_is_result_nan__1_comb = p1_and_7345 | p1_and_7346 | p2_has_0_arg__1_comb & p2_has_inf_arg__1_comb;
  assign p2_is_result_nan__2_comb = p1_and_7343 | p1_and_7344 | p2_has_0_arg__2_comb & p2_has_inf_arg__2_comb;
  assign p2_is_result_nan__4_comb = p1_and_7345 | p1_and_7344 | p2_has_0_arg__4_comb & p2_has_inf_arg__4_comb;
  assign p2_is_result_nan__3_comb = p1_and_7343 | p1_and_7346 | p2_has_0_arg__3_comb & p2_has_inf_arg__3_comb;
  assign p2_fraction__2_comb = p2_fraction__1_comb >> p2_fraction__1_comb[47];
  assign p2_sticky__1_comb = {47'h0000_0000_0000, p2_fraction__1_comb[0]};
  assign p2_fraction__9_comb = p2_fraction__8_comb >> p2_fraction__8_comb[47];
  assign p2_sticky__2_comb = {47'h0000_0000_0000, p2_fraction__8_comb[0]};
  assign p2_fraction__17_comb = p2_fraction__16_comb >> p2_fraction__16_comb[47];
  assign p2_sticky__4_comb = {47'h0000_0000_0000, p2_fraction__16_comb[0]};
  assign p2_fraction__25_comb = p2_fraction__24_comb >> p2_fraction__24_comb[47];
  assign p2_sticky__6_comb = {47'h0000_0000_0000, p2_fraction__24_comb[0]};
  assign p2_exp__2_comb = p2_exp__1_comb & {10{~(p1_eq_7308 | p1_eq_7309)}};
  assign p2_exp__5_comb = p2_exp__4_comb & {10{~(p1_eq_7311 | p1_eq_7312)}};
  assign p2_exp__9_comb = p2_exp__8_comb & {10{~(p1_eq_7308 | p1_eq_7312)}};
  assign p2_exp__13_comb = p2_exp__12_comb & {10{~(p1_eq_7311 | p1_eq_7309)}};
  assign p2_fraction__3_comb = p2_fraction__2_comb | p2_sticky__1_comb;
  assign p2_fraction__10_comb = p2_fraction__9_comb | p2_sticky__2_comb;
  assign p2_fraction__18_comb = p2_fraction__17_comb | p2_sticky__4_comb;
  assign p2_fraction__26_comb = p2_fraction__25_comb | p2_sticky__6_comb;
  assign p2_exp__3_comb = p2_exp__2_comb + {9'h000, p2_fraction__1_comb[47]};
  assign p2_exp__6_comb = p2_exp__5_comb + {9'h000, p2_fraction__8_comb[47]};
  assign p2_exp__10_comb = p2_exp__9_comb + {9'h000, p2_fraction__16_comb[47]};
  assign p2_exp__14_comb = p2_exp__13_comb + {9'h000, p2_fraction__24_comb[47]};
  assign p2_nor_7497_comb = ~(p1_and_7333 | p1_and_7334);
  assign p2_nor_7499_comb = ~(p1_and_7337 | p1_and_7338);
  assign p2_nor_7501_comb = ~(p1_and_7333 | p1_and_7338);
  assign p2_nor_7503_comb = ~(p1_and_7337 | p1_and_7334);
  assign p2_result_sign__3_comb = ~p2_is_result_nan__1_comb & p1_result_sign__2;
  assign p2_result_sign__5_comb = ~p2_is_result_nan__2_comb & p1_result_sign__1;
  assign p2_result_sign__8_comb = ~p2_is_result_nan__4_comb & p1_result_sign__6;
  assign p2_result_sign__7_comb = ~p2_is_result_nan__3_comb & p1_result_sign__4;

  // Registers for pipe stage 2:
  reg [47:0] p2_fraction__3;
  reg [47:0] p2_fraction__10;
  reg [47:0] p2_fraction__18;
  reg [47:0] p2_fraction__26;
  reg [9:0] p2_exp__3;
  reg [9:0] p2_exp__6;
  reg [9:0] p2_exp__10;
  reg [9:0] p2_exp__14;
  reg p2_has_inf_arg__2;
  reg p2_has_inf_arg__1;
  reg p2_has_inf_arg__3;
  reg p2_has_inf_arg__4;
  reg p2_nor_7497;
  reg p2_nor_7499;
  reg p2_nor_7501;
  reg p2_nor_7503;
  reg p2_is_result_nan__2;
  reg p2_is_result_nan__1;
  reg p2_is_result_nan__3;
  reg p2_is_result_nan__4;
  reg p2_result_sign__3;
  reg p2_result_sign__5;
  reg p2_result_sign__8;
  reg p2_result_sign__7;
  reg [22:0] p2_in0_r_fraction__6;
  reg [7:0] p2_in0_r_bexp__6;
  reg [22:0] p2_in0_i_fraction__6;
  reg [7:0] p2_in0_i_bexp__6;
  reg p2_in0_r_sign__2;
  reg p2_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p2_fraction__3 <= p2_fraction__3_comb;
    p2_fraction__10 <= p2_fraction__10_comb;
    p2_fraction__18 <= p2_fraction__18_comb;
    p2_fraction__26 <= p2_fraction__26_comb;
    p2_exp__3 <= p2_exp__3_comb;
    p2_exp__6 <= p2_exp__6_comb;
    p2_exp__10 <= p2_exp__10_comb;
    p2_exp__14 <= p2_exp__14_comb;
    p2_has_inf_arg__2 <= p2_has_inf_arg__2_comb;
    p2_has_inf_arg__1 <= p2_has_inf_arg__1_comb;
    p2_has_inf_arg__3 <= p2_has_inf_arg__3_comb;
    p2_has_inf_arg__4 <= p2_has_inf_arg__4_comb;
    p2_nor_7497 <= p2_nor_7497_comb;
    p2_nor_7499 <= p2_nor_7499_comb;
    p2_nor_7501 <= p2_nor_7501_comb;
    p2_nor_7503 <= p2_nor_7503_comb;
    p2_is_result_nan__2 <= p2_is_result_nan__2_comb;
    p2_is_result_nan__1 <= p2_is_result_nan__1_comb;
    p2_is_result_nan__3 <= p2_is_result_nan__3_comb;
    p2_is_result_nan__4 <= p2_is_result_nan__4_comb;
    p2_result_sign__3 <= p2_result_sign__3_comb;
    p2_result_sign__5 <= p2_result_sign__5_comb;
    p2_result_sign__8 <= p2_result_sign__8_comb;
    p2_result_sign__7 <= p2_result_sign__7_comb;
    p2_in0_r_fraction__6 <= p1_in0_r_fraction__6;
    p2_in0_r_bexp__6 <= p1_in0_r_bexp__6;
    p2_in0_i_fraction__6 <= p1_in0_i_fraction__6;
    p2_in0_i_bexp__6 <= p1_in0_i_bexp__6;
    p2_in0_r_sign__2 <= p1_in0_r_sign__2;
    p2_in0_i_sign__2 <= p1_in0_i_sign__2;
  end

  // ===== Pipe stage 3:
  wire [47:0] p3_fraction__4_comb;
  wire [47:0] p3_sticky__5_comb;
  wire [47:0] p3_fraction__11_comb;
  wire [47:0] p3_sticky__3_comb;
  wire [47:0] p3_fraction__19_comb;
  wire [47:0] p3_sticky__7_comb;
  wire [47:0] p3_fraction__27_comb;
  wire [47:0] p3_sticky__8_comb;
  wire [47:0] p3_fraction__5_comb;
  wire [47:0] p3_fraction__12_comb;
  wire [47:0] p3_fraction__20_comb;
  wire [47:0] p3_fraction__28_comb;
  wire [21:0] p3_bit_slice_7617_comb;
  wire [21:0] p3_bit_slice_7618_comb;
  wire [21:0] p3_bit_slice_7619_comb;
  wire [21:0] p3_bit_slice_7620_comb;
  wire p3_bit_slice_7621_comb;
  wire p3_bit_slice_7622_comb;
  wire [22:0] p3_fraction__6_comb;
  wire p3_bit_slice_7624_comb;
  wire p3_bit_slice_7625_comb;
  wire [22:0] p3_fraction__13_comb;
  wire p3_bit_slice_7627_comb;
  wire p3_bit_slice_7628_comb;
  wire [22:0] p3_fraction__21_comb;
  wire p3_bit_slice_7630_comb;
  wire p3_bit_slice_7631_comb;
  wire [22:0] p3_fraction__29_comb;
  wire p3_bd__1_sign_comb;
  assign p3_fraction__4_comb = $signed(p2_exp__3) <= $signed(10'h000) ? {1'h0, p2_fraction__3[47:1]} : p2_fraction__3;
  assign p3_sticky__5_comb = {47'h0000_0000_0000, p2_fraction__3[0]};
  assign p3_fraction__11_comb = $signed(p2_exp__6) <= $signed(10'h000) ? {1'h0, p2_fraction__10[47:1]} : p2_fraction__10;
  assign p3_sticky__3_comb = {47'h0000_0000_0000, p2_fraction__10[0]};
  assign p3_fraction__19_comb = $signed(p2_exp__10) <= $signed(10'h000) ? {1'h0, p2_fraction__18[47:1]} : p2_fraction__18;
  assign p3_sticky__7_comb = {47'h0000_0000_0000, p2_fraction__18[0]};
  assign p3_fraction__27_comb = $signed(p2_exp__14) <= $signed(10'h000) ? {1'h0, p2_fraction__26[47:1]} : p2_fraction__26;
  assign p3_sticky__8_comb = {47'h0000_0000_0000, p2_fraction__26[0]};
  assign p3_fraction__5_comb = p3_fraction__4_comb | p3_sticky__5_comb;
  assign p3_fraction__12_comb = p3_fraction__11_comb | p3_sticky__3_comb;
  assign p3_fraction__20_comb = p3_fraction__19_comb | p3_sticky__7_comb;
  assign p3_fraction__28_comb = p3_fraction__27_comb | p3_sticky__8_comb;
  assign p3_bit_slice_7617_comb = p3_fraction__5_comb[21:0];
  assign p3_bit_slice_7618_comb = p3_fraction__12_comb[21:0];
  assign p3_bit_slice_7619_comb = p3_fraction__20_comb[21:0];
  assign p3_bit_slice_7620_comb = p3_fraction__28_comb[21:0];
  assign p3_bit_slice_7621_comb = p3_fraction__5_comb[22];
  assign p3_bit_slice_7622_comb = p3_fraction__5_comb[23];
  assign p3_fraction__6_comb = p3_fraction__5_comb[45:23];
  assign p3_bit_slice_7624_comb = p3_fraction__12_comb[22];
  assign p3_bit_slice_7625_comb = p3_fraction__12_comb[23];
  assign p3_fraction__13_comb = p3_fraction__12_comb[45:23];
  assign p3_bit_slice_7627_comb = p3_fraction__20_comb[22];
  assign p3_bit_slice_7628_comb = p3_fraction__20_comb[23];
  assign p3_fraction__21_comb = p3_fraction__20_comb[45:23];
  assign p3_bit_slice_7630_comb = p3_fraction__28_comb[22];
  assign p3_bit_slice_7631_comb = p3_fraction__28_comb[23];
  assign p3_fraction__29_comb = p3_fraction__28_comb[45:23];
  assign p3_bd__1_sign_comb = ~p2_result_sign__3;

  // Registers for pipe stage 3:
  reg [9:0] p3_exp__3;
  reg [9:0] p3_exp__6;
  reg [9:0] p3_exp__10;
  reg [9:0] p3_exp__14;
  reg [21:0] p3_bit_slice_7617;
  reg [21:0] p3_bit_slice_7618;
  reg [21:0] p3_bit_slice_7619;
  reg [21:0] p3_bit_slice_7620;
  reg p3_bit_slice_7621;
  reg p3_bit_slice_7622;
  reg [22:0] p3_fraction__6;
  reg p3_bit_slice_7624;
  reg p3_bit_slice_7625;
  reg [22:0] p3_fraction__13;
  reg p3_bit_slice_7627;
  reg p3_bit_slice_7628;
  reg [22:0] p3_fraction__21;
  reg p3_bit_slice_7630;
  reg p3_bit_slice_7631;
  reg [22:0] p3_fraction__29;
  reg p3_has_inf_arg__2;
  reg p3_has_inf_arg__1;
  reg p3_has_inf_arg__3;
  reg p3_has_inf_arg__4;
  reg p3_nor_7497;
  reg p3_nor_7499;
  reg p3_nor_7501;
  reg p3_nor_7503;
  reg p3_is_result_nan__2;
  reg p3_is_result_nan__1;
  reg p3_is_result_nan__3;
  reg p3_is_result_nan__4;
  reg p3_bd__1_sign;
  reg p3_result_sign__5;
  reg p3_result_sign__8;
  reg p3_result_sign__7;
  reg [22:0] p3_in0_r_fraction__6;
  reg [7:0] p3_in0_r_bexp__6;
  reg [22:0] p3_in0_i_fraction__6;
  reg [7:0] p3_in0_i_bexp__6;
  reg p3_in0_r_sign__2;
  reg p3_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p3_exp__3 <= p2_exp__3;
    p3_exp__6 <= p2_exp__6;
    p3_exp__10 <= p2_exp__10;
    p3_exp__14 <= p2_exp__14;
    p3_bit_slice_7617 <= p3_bit_slice_7617_comb;
    p3_bit_slice_7618 <= p3_bit_slice_7618_comb;
    p3_bit_slice_7619 <= p3_bit_slice_7619_comb;
    p3_bit_slice_7620 <= p3_bit_slice_7620_comb;
    p3_bit_slice_7621 <= p3_bit_slice_7621_comb;
    p3_bit_slice_7622 <= p3_bit_slice_7622_comb;
    p3_fraction__6 <= p3_fraction__6_comb;
    p3_bit_slice_7624 <= p3_bit_slice_7624_comb;
    p3_bit_slice_7625 <= p3_bit_slice_7625_comb;
    p3_fraction__13 <= p3_fraction__13_comb;
    p3_bit_slice_7627 <= p3_bit_slice_7627_comb;
    p3_bit_slice_7628 <= p3_bit_slice_7628_comb;
    p3_fraction__21 <= p3_fraction__21_comb;
    p3_bit_slice_7630 <= p3_bit_slice_7630_comb;
    p3_bit_slice_7631 <= p3_bit_slice_7631_comb;
    p3_fraction__29 <= p3_fraction__29_comb;
    p3_has_inf_arg__2 <= p2_has_inf_arg__2;
    p3_has_inf_arg__1 <= p2_has_inf_arg__1;
    p3_has_inf_arg__3 <= p2_has_inf_arg__3;
    p3_has_inf_arg__4 <= p2_has_inf_arg__4;
    p3_nor_7497 <= p2_nor_7497;
    p3_nor_7499 <= p2_nor_7499;
    p3_nor_7501 <= p2_nor_7501;
    p3_nor_7503 <= p2_nor_7503;
    p3_is_result_nan__2 <= p2_is_result_nan__2;
    p3_is_result_nan__1 <= p2_is_result_nan__1;
    p3_is_result_nan__3 <= p2_is_result_nan__3;
    p3_is_result_nan__4 <= p2_is_result_nan__4;
    p3_bd__1_sign <= p3_bd__1_sign_comb;
    p3_result_sign__5 <= p2_result_sign__5;
    p3_result_sign__8 <= p2_result_sign__8;
    p3_result_sign__7 <= p2_result_sign__7;
    p3_in0_r_fraction__6 <= p2_in0_r_fraction__6;
    p3_in0_r_bexp__6 <= p2_in0_r_bexp__6;
    p3_in0_i_fraction__6 <= p2_in0_i_fraction__6;
    p3_in0_i_bexp__6 <= p2_in0_i_bexp__6;
    p3_in0_r_sign__2 <= p2_in0_r_sign__2;
    p3_in0_i_sign__2 <= p2_in0_i_sign__2;
  end

  // ===== Pipe stage 4:
  wire p4_greater_than_half_way__2_comb;
  wire [23:0] p4_fraction__7_comb;
  wire p4_greater_than_half_way__1_comb;
  wire [23:0] p4_fraction__14_comb;
  wire p4_greater_than_half_way__3_comb;
  wire [23:0] p4_fraction__22_comb;
  wire p4_greater_than_half_way__4_comb;
  wire [23:0] p4_fraction__30_comb;
  wire p4_do_round_up__2_comb;
  wire [23:0] p4_add_7755_comb;
  wire p4_do_round_up__1_comb;
  wire [23:0] p4_add_7757_comb;
  wire p4_do_round_up__3_comb;
  wire [23:0] p4_add_7759_comb;
  wire p4_do_round_up__4_comb;
  wire [23:0] p4_add_7761_comb;
  wire [23:0] p4_fraction__23_comb;
  wire [23:0] p4_fraction__15_comb;
  wire [23:0] p4_fraction__31_comb;
  wire [23:0] p4_fraction__32_comb;
  assign p4_greater_than_half_way__2_comb = p3_bit_slice_7621 & p3_bit_slice_7617 != 22'h00_0000;
  assign p4_fraction__7_comb = {1'h0, p3_fraction__6};
  assign p4_greater_than_half_way__1_comb = p3_bit_slice_7624 & p3_bit_slice_7618 != 22'h00_0000;
  assign p4_fraction__14_comb = {1'h0, p3_fraction__13};
  assign p4_greater_than_half_way__3_comb = p3_bit_slice_7627 & p3_bit_slice_7619 != 22'h00_0000;
  assign p4_fraction__22_comb = {1'h0, p3_fraction__21};
  assign p4_greater_than_half_way__4_comb = p3_bit_slice_7630 & p3_bit_slice_7620 != 22'h00_0000;
  assign p4_fraction__30_comb = {1'h0, p3_fraction__29};
  assign p4_do_round_up__2_comb = p4_greater_than_half_way__2_comb | p3_bit_slice_7621 & p3_bit_slice_7617 == 22'h00_0000 & p3_bit_slice_7622;
  assign p4_add_7755_comb = p4_fraction__7_comb + 24'h00_0001;
  assign p4_do_round_up__1_comb = p4_greater_than_half_way__1_comb | p3_bit_slice_7624 & p3_bit_slice_7618 == 22'h00_0000 & p3_bit_slice_7625;
  assign p4_add_7757_comb = p4_fraction__14_comb + 24'h00_0001;
  assign p4_do_round_up__3_comb = p4_greater_than_half_way__3_comb | p3_bit_slice_7627 & p3_bit_slice_7619 == 22'h00_0000 & p3_bit_slice_7628;
  assign p4_add_7759_comb = p4_fraction__22_comb + 24'h00_0001;
  assign p4_do_round_up__4_comb = p4_greater_than_half_way__4_comb | p3_bit_slice_7630 & p3_bit_slice_7620 == 22'h00_0000 & p3_bit_slice_7631;
  assign p4_add_7761_comb = p4_fraction__30_comb + 24'h00_0001;
  assign p4_fraction__23_comb = p4_do_round_up__2_comb ? p4_add_7755_comb : p4_fraction__7_comb;
  assign p4_fraction__15_comb = p4_do_round_up__1_comb ? p4_add_7757_comb : p4_fraction__14_comb;
  assign p4_fraction__31_comb = p4_do_round_up__3_comb ? p4_add_7759_comb : p4_fraction__22_comb;
  assign p4_fraction__32_comb = p4_do_round_up__4_comb ? p4_add_7761_comb : p4_fraction__30_comb;

  // Registers for pipe stage 4:
  reg [9:0] p4_exp__3;
  reg [9:0] p4_exp__6;
  reg [9:0] p4_exp__10;
  reg [9:0] p4_exp__14;
  reg [23:0] p4_fraction__23;
  reg [23:0] p4_fraction__15;
  reg [23:0] p4_fraction__31;
  reg [23:0] p4_fraction__32;
  reg p4_has_inf_arg__2;
  reg p4_has_inf_arg__1;
  reg p4_has_inf_arg__3;
  reg p4_has_inf_arg__4;
  reg p4_nor_7497;
  reg p4_nor_7499;
  reg p4_nor_7501;
  reg p4_nor_7503;
  reg p4_is_result_nan__2;
  reg p4_is_result_nan__1;
  reg p4_is_result_nan__3;
  reg p4_is_result_nan__4;
  reg p4_bd__1_sign;
  reg p4_result_sign__5;
  reg p4_result_sign__8;
  reg p4_result_sign__7;
  reg [22:0] p4_in0_r_fraction__6;
  reg [7:0] p4_in0_r_bexp__6;
  reg [22:0] p4_in0_i_fraction__6;
  reg [7:0] p4_in0_i_bexp__6;
  reg p4_in0_r_sign__2;
  reg p4_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p4_exp__3 <= p3_exp__3;
    p4_exp__6 <= p3_exp__6;
    p4_exp__10 <= p3_exp__10;
    p4_exp__14 <= p3_exp__14;
    p4_fraction__23 <= p4_fraction__23_comb;
    p4_fraction__15 <= p4_fraction__15_comb;
    p4_fraction__31 <= p4_fraction__31_comb;
    p4_fraction__32 <= p4_fraction__32_comb;
    p4_has_inf_arg__2 <= p3_has_inf_arg__2;
    p4_has_inf_arg__1 <= p3_has_inf_arg__1;
    p4_has_inf_arg__3 <= p3_has_inf_arg__3;
    p4_has_inf_arg__4 <= p3_has_inf_arg__4;
    p4_nor_7497 <= p3_nor_7497;
    p4_nor_7499 <= p3_nor_7499;
    p4_nor_7501 <= p3_nor_7501;
    p4_nor_7503 <= p3_nor_7503;
    p4_is_result_nan__2 <= p3_is_result_nan__2;
    p4_is_result_nan__1 <= p3_is_result_nan__1;
    p4_is_result_nan__3 <= p3_is_result_nan__3;
    p4_is_result_nan__4 <= p3_is_result_nan__4;
    p4_bd__1_sign <= p3_bd__1_sign;
    p4_result_sign__5 <= p3_result_sign__5;
    p4_result_sign__8 <= p3_result_sign__8;
    p4_result_sign__7 <= p3_result_sign__7;
    p4_in0_r_fraction__6 <= p3_in0_r_fraction__6;
    p4_in0_r_bexp__6 <= p3_in0_r_bexp__6;
    p4_in0_i_fraction__6 <= p3_in0_i_fraction__6;
    p4_in0_i_bexp__6 <= p3_in0_i_bexp__6;
    p4_in0_r_sign__2 <= p3_in0_r_sign__2;
    p4_in0_i_sign__2 <= p3_in0_i_sign__2;
  end

  // ===== Pipe stage 5:
  wire [9:0] p5_add_7831_comb;
  wire [9:0] p5_add_7833_comb;
  wire [9:0] p5_add_7835_comb;
  wire [9:0] p5_add_7837_comb;
  wire [9:0] p5_exp__11_comb;
  wire [9:0] p5_exp__7_comb;
  wire [9:0] p5_exp__15_comb;
  wire [9:0] p5_exp__16_comb;
  wire p5_sgt_7846_comb;
  wire p5_sgt_7847_comb;
  wire p5_sgt_7848_comb;
  wire p5_sgt_7849_comb;
  wire [8:0] p5_result_exp__1_comb;
  wire [8:0] p5_result_exp__2_comb;
  wire [8:0] p5_result_exp__6_comb;
  wire [8:0] p5_result_exp__9_comb;
  wire [22:0] p5_result_fraction__3_comb;
  wire [22:0] p5_result_fraction__1_comb;
  wire [22:0] p5_result_fraction__6_comb;
  wire [22:0] p5_result_fraction__9_comb;
  assign p5_add_7831_comb = p4_exp__3 + 10'h001;
  assign p5_add_7833_comb = p4_exp__6 + 10'h001;
  assign p5_add_7835_comb = p4_exp__10 + 10'h001;
  assign p5_add_7837_comb = p4_exp__14 + 10'h001;
  assign p5_exp__11_comb = p4_fraction__23[23] ? p5_add_7831_comb : p4_exp__3;
  assign p5_exp__7_comb = p4_fraction__15[23] ? p5_add_7833_comb : p4_exp__6;
  assign p5_exp__15_comb = p4_fraction__31[23] ? p5_add_7835_comb : p4_exp__10;
  assign p5_exp__16_comb = p4_fraction__32[23] ? p5_add_7837_comb : p4_exp__14;
  assign p5_sgt_7846_comb = $signed(p5_exp__11_comb) > $signed(10'h000);
  assign p5_sgt_7847_comb = $signed(p5_exp__7_comb) > $signed(10'h000);
  assign p5_sgt_7848_comb = $signed(p5_exp__15_comb) > $signed(10'h000);
  assign p5_sgt_7849_comb = $signed(p5_exp__16_comb) > $signed(10'h000);
  assign p5_result_exp__1_comb = p5_exp__11_comb[8:0];
  assign p5_result_exp__2_comb = p5_exp__7_comb[8:0];
  assign p5_result_exp__6_comb = p5_exp__15_comb[8:0];
  assign p5_result_exp__9_comb = p5_exp__16_comb[8:0];
  assign p5_result_fraction__3_comb = p4_fraction__23[22:0];
  assign p5_result_fraction__1_comb = p4_fraction__15[22:0];
  assign p5_result_fraction__6_comb = p4_fraction__31[22:0];
  assign p5_result_fraction__9_comb = p4_fraction__32[22:0];

  // Registers for pipe stage 5:
  reg p5_sgt_7846;
  reg p5_sgt_7847;
  reg p5_sgt_7848;
  reg p5_sgt_7849;
  reg [8:0] p5_result_exp__1;
  reg [8:0] p5_result_exp__2;
  reg [8:0] p5_result_exp__6;
  reg [8:0] p5_result_exp__9;
  reg p5_has_inf_arg__2;
  reg p5_has_inf_arg__1;
  reg p5_has_inf_arg__3;
  reg p5_has_inf_arg__4;
  reg p5_nor_7497;
  reg p5_nor_7499;
  reg p5_nor_7501;
  reg p5_nor_7503;
  reg [22:0] p5_result_fraction__3;
  reg p5_is_result_nan__2;
  reg [22:0] p5_result_fraction__1;
  reg p5_is_result_nan__1;
  reg [22:0] p5_result_fraction__6;
  reg p5_is_result_nan__3;
  reg [22:0] p5_result_fraction__9;
  reg p5_is_result_nan__4;
  reg p5_bd__1_sign;
  reg p5_result_sign__5;
  reg p5_result_sign__8;
  reg p5_result_sign__7;
  reg [22:0] p5_in0_r_fraction__6;
  reg [7:0] p5_in0_r_bexp__6;
  reg [22:0] p5_in0_i_fraction__6;
  reg [7:0] p5_in0_i_bexp__6;
  reg p5_in0_r_sign__2;
  reg p5_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p5_sgt_7846 <= p5_sgt_7846_comb;
    p5_sgt_7847 <= p5_sgt_7847_comb;
    p5_sgt_7848 <= p5_sgt_7848_comb;
    p5_sgt_7849 <= p5_sgt_7849_comb;
    p5_result_exp__1 <= p5_result_exp__1_comb;
    p5_result_exp__2 <= p5_result_exp__2_comb;
    p5_result_exp__6 <= p5_result_exp__6_comb;
    p5_result_exp__9 <= p5_result_exp__9_comb;
    p5_has_inf_arg__2 <= p4_has_inf_arg__2;
    p5_has_inf_arg__1 <= p4_has_inf_arg__1;
    p5_has_inf_arg__3 <= p4_has_inf_arg__3;
    p5_has_inf_arg__4 <= p4_has_inf_arg__4;
    p5_nor_7497 <= p4_nor_7497;
    p5_nor_7499 <= p4_nor_7499;
    p5_nor_7501 <= p4_nor_7501;
    p5_nor_7503 <= p4_nor_7503;
    p5_result_fraction__3 <= p5_result_fraction__3_comb;
    p5_is_result_nan__2 <= p4_is_result_nan__2;
    p5_result_fraction__1 <= p5_result_fraction__1_comb;
    p5_is_result_nan__1 <= p4_is_result_nan__1;
    p5_result_fraction__6 <= p5_result_fraction__6_comb;
    p5_is_result_nan__3 <= p4_is_result_nan__3;
    p5_result_fraction__9 <= p5_result_fraction__9_comb;
    p5_is_result_nan__4 <= p4_is_result_nan__4;
    p5_bd__1_sign <= p4_bd__1_sign;
    p5_result_sign__5 <= p4_result_sign__5;
    p5_result_sign__8 <= p4_result_sign__8;
    p5_result_sign__7 <= p4_result_sign__7;
    p5_in0_r_fraction__6 <= p4_in0_r_fraction__6;
    p5_in0_r_bexp__6 <= p4_in0_r_bexp__6;
    p5_in0_i_fraction__6 <= p4_in0_i_fraction__6;
    p5_in0_i_bexp__6 <= p4_in0_i_bexp__6;
    p5_in0_r_sign__2 <= p4_in0_r_sign__2;
    p5_in0_i_sign__2 <= p4_in0_i_sign__2;
  end

  // ===== Pipe stage 6:
  wire [8:0] p6_result_exp__4_comb;
  wire [8:0] p6_result_exp__3_comb;
  wire [8:0] p6_result_exp__7_comb;
  wire [8:0] p6_result_exp__10_comb;
  wire p6_nor_7974_comb;
  wire p6_nor_7975_comb;
  wire p6_nor_7976_comb;
  wire p6_nor_7977_comb;
  wire [7:0] p6_bit_slice_7978_comb;
  wire [7:0] p6_bit_slice_7979_comb;
  wire [7:0] p6_bit_slice_7980_comb;
  wire [7:0] p6_bit_slice_7981_comb;
  assign p6_result_exp__4_comb = p5_result_exp__1 & {9{p5_sgt_7846}};
  assign p6_result_exp__3_comb = p5_result_exp__2 & {9{p5_sgt_7847}};
  assign p6_result_exp__7_comb = p5_result_exp__6 & {9{p5_sgt_7848}};
  assign p6_result_exp__10_comb = p5_result_exp__9 & {9{p5_sgt_7849}};
  assign p6_nor_7974_comb = ~(p6_result_exp__4_comb[8] | p6_result_exp__4_comb[0] & p6_result_exp__4_comb[1] & p6_result_exp__4_comb[2] & p6_result_exp__4_comb[3] & p6_result_exp__4_comb[4] & p6_result_exp__4_comb[5] & p6_result_exp__4_comb[6] & p6_result_exp__4_comb[7]);
  assign p6_nor_7975_comb = ~(p6_result_exp__3_comb[8] | p6_result_exp__3_comb[0] & p6_result_exp__3_comb[1] & p6_result_exp__3_comb[2] & p6_result_exp__3_comb[3] & p6_result_exp__3_comb[4] & p6_result_exp__3_comb[5] & p6_result_exp__3_comb[6] & p6_result_exp__3_comb[7]);
  assign p6_nor_7976_comb = ~(p6_result_exp__7_comb[8] | p6_result_exp__7_comb[0] & p6_result_exp__7_comb[1] & p6_result_exp__7_comb[2] & p6_result_exp__7_comb[3] & p6_result_exp__7_comb[4] & p6_result_exp__7_comb[5] & p6_result_exp__7_comb[6] & p6_result_exp__7_comb[7]);
  assign p6_nor_7977_comb = ~(p6_result_exp__10_comb[8] | p6_result_exp__10_comb[0] & p6_result_exp__10_comb[1] & p6_result_exp__10_comb[2] & p6_result_exp__10_comb[3] & p6_result_exp__10_comb[4] & p6_result_exp__10_comb[5] & p6_result_exp__10_comb[6] & p6_result_exp__10_comb[7]);
  assign p6_bit_slice_7978_comb = p6_result_exp__4_comb[7:0];
  assign p6_bit_slice_7979_comb = p6_result_exp__3_comb[7:0];
  assign p6_bit_slice_7980_comb = p6_result_exp__7_comb[7:0];
  assign p6_bit_slice_7981_comb = p6_result_exp__10_comb[7:0];

  // Registers for pipe stage 6:
  reg p6_sgt_7846;
  reg p6_sgt_7847;
  reg p6_sgt_7848;
  reg p6_sgt_7849;
  reg p6_has_inf_arg__2;
  reg p6_has_inf_arg__1;
  reg p6_has_inf_arg__3;
  reg p6_has_inf_arg__4;
  reg p6_nor_7974;
  reg p6_nor_7497;
  reg p6_nor_7975;
  reg p6_nor_7499;
  reg p6_nor_7976;
  reg p6_nor_7501;
  reg p6_nor_7977;
  reg p6_nor_7503;
  reg [22:0] p6_result_fraction__3;
  reg p6_is_result_nan__2;
  reg [22:0] p6_result_fraction__1;
  reg p6_is_result_nan__1;
  reg [22:0] p6_result_fraction__6;
  reg p6_is_result_nan__3;
  reg [22:0] p6_result_fraction__9;
  reg p6_is_result_nan__4;
  reg [7:0] p6_bit_slice_7978;
  reg [7:0] p6_bit_slice_7979;
  reg [7:0] p6_bit_slice_7980;
  reg [7:0] p6_bit_slice_7981;
  reg p6_bd__1_sign;
  reg p6_result_sign__5;
  reg p6_result_sign__8;
  reg p6_result_sign__7;
  reg [22:0] p6_in0_r_fraction__6;
  reg [7:0] p6_in0_r_bexp__6;
  reg [22:0] p6_in0_i_fraction__6;
  reg [7:0] p6_in0_i_bexp__6;
  reg p6_in0_r_sign__2;
  reg p6_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p6_sgt_7846 <= p5_sgt_7846;
    p6_sgt_7847 <= p5_sgt_7847;
    p6_sgt_7848 <= p5_sgt_7848;
    p6_sgt_7849 <= p5_sgt_7849;
    p6_has_inf_arg__2 <= p5_has_inf_arg__2;
    p6_has_inf_arg__1 <= p5_has_inf_arg__1;
    p6_has_inf_arg__3 <= p5_has_inf_arg__3;
    p6_has_inf_arg__4 <= p5_has_inf_arg__4;
    p6_nor_7974 <= p6_nor_7974_comb;
    p6_nor_7497 <= p5_nor_7497;
    p6_nor_7975 <= p6_nor_7975_comb;
    p6_nor_7499 <= p5_nor_7499;
    p6_nor_7976 <= p6_nor_7976_comb;
    p6_nor_7501 <= p5_nor_7501;
    p6_nor_7977 <= p6_nor_7977_comb;
    p6_nor_7503 <= p5_nor_7503;
    p6_result_fraction__3 <= p5_result_fraction__3;
    p6_is_result_nan__2 <= p5_is_result_nan__2;
    p6_result_fraction__1 <= p5_result_fraction__1;
    p6_is_result_nan__1 <= p5_is_result_nan__1;
    p6_result_fraction__6 <= p5_result_fraction__6;
    p6_is_result_nan__3 <= p5_is_result_nan__3;
    p6_result_fraction__9 <= p5_result_fraction__9;
    p6_is_result_nan__4 <= p5_is_result_nan__4;
    p6_bit_slice_7978 <= p6_bit_slice_7978_comb;
    p6_bit_slice_7979 <= p6_bit_slice_7979_comb;
    p6_bit_slice_7980 <= p6_bit_slice_7980_comb;
    p6_bit_slice_7981 <= p6_bit_slice_7981_comb;
    p6_bd__1_sign <= p5_bd__1_sign;
    p6_result_sign__5 <= p5_result_sign__5;
    p6_result_sign__8 <= p5_result_sign__8;
    p6_result_sign__7 <= p5_result_sign__7;
    p6_in0_r_fraction__6 <= p5_in0_r_fraction__6;
    p6_in0_r_bexp__6 <= p5_in0_r_bexp__6;
    p6_in0_i_fraction__6 <= p5_in0_i_fraction__6;
    p6_in0_i_bexp__6 <= p5_in0_i_bexp__6;
    p6_in0_r_sign__2 <= p5_in0_r_sign__2;
    p6_in0_i_sign__2 <= p5_in0_i_sign__2;
  end

  // ===== Pipe stage 7:
  wire [22:0] p7_result_fraction__4_comb;
  wire [22:0] p7_nan_fraction__1_comb;
  wire [7:0] p7_high_exp__29_comb;
  wire [22:0] p7_result_fraction__2_comb;
  wire [22:0] p7_nan_fraction__5_comb;
  wire [7:0] p7_high_exp__28_comb;
  wire [22:0] p7_result_fraction__7_comb;
  wire [22:0] p7_nan_fraction__3_comb;
  wire [7:0] p7_high_exp__30_comb;
  wire [22:0] p7_result_fraction__10_comb;
  wire [22:0] p7_nan_fraction__4_comb;
  wire [7:0] p7_high_exp__31_comb;
  wire [22:0] p7_result_fraction__8_comb;
  wire [7:0] p7_result_exp__8_comb;
  wire [22:0] p7_result_fraction__5_comb;
  wire [7:0] p7_result_exp__5_comb;
  wire [22:0] p7_result_fraction__11_comb;
  wire [7:0] p7_result_exp__11_comb;
  wire [22:0] p7_result_fraction__12_comb;
  wire [7:0] p7_result_exp__12_comb;
  wire [24:0] p7_or_8122_comb;
  wire p7_ne_8124_comb;
  wire [5:0] p7_add_8125_comb;
  wire [1:0] p7_bit_slice_8126_comb;
  wire p7_ugt_8127_comb;
  wire [24:0] p7_or_8128_comb;
  wire p7_ne_8130_comb;
  wire [5:0] p7_add_8131_comb;
  wire [1:0] p7_bit_slice_8132_comb;
  wire [24:0] p7_or_8133_comb;
  wire p7_ne_8135_comb;
  wire [5:0] p7_add_8136_comb;
  wire [1:0] p7_bit_slice_8137_comb;
  wire p7_ugt_8138_comb;
  wire [24:0] p7_or_8139_comb;
  wire p7_ne_8141_comb;
  wire [5:0] p7_add_8142_comb;
  wire [1:0] p7_bit_slice_8143_comb;
  wire p7_eq_8148_comb;
  wire p7_eq_8149_comb;
  wire p7_eq_8150_comb;
  wire p7_eq_8151_comb;
  wire p7_ne_8156_comb;
  wire p7_ne_8157_comb;
  wire p7_ne_8158_comb;
  wire p7_ne_8159_comb;
  assign p7_result_fraction__4_comb = p6_result_fraction__3 & {23{p6_sgt_7846}} & {23{p6_nor_7974}} & {23{p6_nor_7497}};
  assign p7_nan_fraction__1_comb = 23'h40_0000;
  assign p7_high_exp__29_comb = 8'hff;
  assign p7_result_fraction__2_comb = p6_result_fraction__1 & {23{p6_sgt_7847}} & {23{p6_nor_7975}} & {23{p6_nor_7499}};
  assign p7_nan_fraction__5_comb = 23'h40_0000;
  assign p7_high_exp__28_comb = 8'hff;
  assign p7_result_fraction__7_comb = p6_result_fraction__6 & {23{p6_sgt_7848}} & {23{p6_nor_7976}} & {23{p6_nor_7501}};
  assign p7_nan_fraction__3_comb = 23'h40_0000;
  assign p7_high_exp__30_comb = 8'hff;
  assign p7_result_fraction__10_comb = p6_result_fraction__9 & {23{p6_sgt_7849}} & {23{p6_nor_7977}} & {23{p6_nor_7503}};
  assign p7_nan_fraction__4_comb = 23'h40_0000;
  assign p7_high_exp__31_comb = 8'hff;
  assign p7_result_fraction__8_comb = p6_is_result_nan__2 ? p7_nan_fraction__1_comb : p7_result_fraction__4_comb;
  assign p7_result_exp__8_comb = p6_is_result_nan__2 | p6_has_inf_arg__2 | ~p6_nor_7974 ? p7_high_exp__29_comb : p6_bit_slice_7978;
  assign p7_result_fraction__5_comb = p6_is_result_nan__1 ? p7_nan_fraction__5_comb : p7_result_fraction__2_comb;
  assign p7_result_exp__5_comb = p6_is_result_nan__1 | p6_has_inf_arg__1 | ~p6_nor_7975 ? p7_high_exp__28_comb : p6_bit_slice_7979;
  assign p7_result_fraction__11_comb = p6_is_result_nan__3 ? p7_nan_fraction__3_comb : p7_result_fraction__7_comb;
  assign p7_result_exp__11_comb = p6_is_result_nan__3 | p6_has_inf_arg__3 | ~p6_nor_7976 ? p7_high_exp__30_comb : p6_bit_slice_7980;
  assign p7_result_fraction__12_comb = p6_is_result_nan__4 ? p7_nan_fraction__4_comb : p7_result_fraction__10_comb;
  assign p7_result_exp__12_comb = p6_is_result_nan__4 | p6_has_inf_arg__4 | ~p6_nor_7977 ? p7_high_exp__31_comb : p6_bit_slice_7981;
  assign p7_or_8122_comb = {2'h0, p7_result_fraction__8_comb} | 25'h080_0000;
  assign p7_ne_8124_comb = p7_result_exp__8_comb != 8'h00;
  assign p7_add_8125_comb = p7_result_exp__8_comb[7:2] + 6'h07;
  assign p7_bit_slice_8126_comb = p7_result_exp__8_comb[1:0];
  assign p7_ugt_8127_comb = p7_result_exp__8_comb > p7_result_exp__5_comb;
  assign p7_or_8128_comb = {2'h0, p7_result_fraction__5_comb} | 25'h080_0000;
  assign p7_ne_8130_comb = p7_result_exp__5_comb != 8'h00;
  assign p7_add_8131_comb = p7_result_exp__5_comb[7:2] + 6'h07;
  assign p7_bit_slice_8132_comb = p7_result_exp__5_comb[1:0];
  assign p7_or_8133_comb = {2'h0, p7_result_fraction__11_comb} | 25'h080_0000;
  assign p7_ne_8135_comb = p7_result_exp__11_comb != 8'h00;
  assign p7_add_8136_comb = p7_result_exp__11_comb[7:2] + 6'h07;
  assign p7_bit_slice_8137_comb = p7_result_exp__11_comb[1:0];
  assign p7_ugt_8138_comb = p7_result_exp__11_comb > p7_result_exp__12_comb;
  assign p7_or_8139_comb = {2'h0, p7_result_fraction__12_comb} | 25'h080_0000;
  assign p7_ne_8141_comb = p7_result_exp__12_comb != 8'h00;
  assign p7_add_8142_comb = p7_result_exp__12_comb[7:2] + 6'h07;
  assign p7_bit_slice_8143_comb = p7_result_exp__12_comb[1:0];
  assign p7_eq_8148_comb = p7_result_fraction__8_comb == 23'h00_0000;
  assign p7_eq_8149_comb = p7_result_fraction__5_comb == 23'h00_0000;
  assign p7_eq_8150_comb = p7_result_fraction__11_comb == 23'h00_0000;
  assign p7_eq_8151_comb = p7_result_fraction__12_comb == 23'h00_0000;
  assign p7_ne_8156_comb = p7_result_fraction__8_comb != 23'h00_0000;
  assign p7_ne_8157_comb = p7_result_fraction__5_comb != 23'h00_0000;
  assign p7_ne_8158_comb = p7_result_fraction__11_comb != 23'h00_0000;
  assign p7_ne_8159_comb = p7_result_fraction__12_comb != 23'h00_0000;

  // Registers for pipe stage 7:
  reg [7:0] p7_result_exp__8;
  reg [7:0] p7_result_exp__5;
  reg [7:0] p7_result_exp__11;
  reg [7:0] p7_result_exp__12;
  reg [24:0] p7_or_8122;
  reg p7_ne_8124;
  reg [5:0] p7_add_8125;
  reg [1:0] p7_bit_slice_8126;
  reg p7_ugt_8127;
  reg [24:0] p7_or_8128;
  reg p7_ne_8130;
  reg [5:0] p7_add_8131;
  reg [1:0] p7_bit_slice_8132;
  reg [24:0] p7_or_8133;
  reg p7_ne_8135;
  reg [5:0] p7_add_8136;
  reg [1:0] p7_bit_slice_8137;
  reg p7_ugt_8138;
  reg [24:0] p7_or_8139;
  reg p7_ne_8141;
  reg [5:0] p7_add_8142;
  reg [1:0] p7_bit_slice_8143;
  reg p7_bd__1_sign;
  reg p7_result_sign__5;
  reg p7_result_sign__8;
  reg p7_result_sign__7;
  reg p7_eq_8148;
  reg p7_eq_8149;
  reg p7_eq_8150;
  reg p7_eq_8151;
  reg p7_ne_8156;
  reg p7_ne_8157;
  reg p7_ne_8158;
  reg p7_ne_8159;
  reg [22:0] p7_in0_r_fraction__6;
  reg [7:0] p7_in0_r_bexp__6;
  reg [22:0] p7_in0_i_fraction__6;
  reg [7:0] p7_in0_i_bexp__6;
  reg p7_in0_r_sign__2;
  reg p7_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p7_result_exp__8 <= p7_result_exp__8_comb;
    p7_result_exp__5 <= p7_result_exp__5_comb;
    p7_result_exp__11 <= p7_result_exp__11_comb;
    p7_result_exp__12 <= p7_result_exp__12_comb;
    p7_or_8122 <= p7_or_8122_comb;
    p7_ne_8124 <= p7_ne_8124_comb;
    p7_add_8125 <= p7_add_8125_comb;
    p7_bit_slice_8126 <= p7_bit_slice_8126_comb;
    p7_ugt_8127 <= p7_ugt_8127_comb;
    p7_or_8128 <= p7_or_8128_comb;
    p7_ne_8130 <= p7_ne_8130_comb;
    p7_add_8131 <= p7_add_8131_comb;
    p7_bit_slice_8132 <= p7_bit_slice_8132_comb;
    p7_or_8133 <= p7_or_8133_comb;
    p7_ne_8135 <= p7_ne_8135_comb;
    p7_add_8136 <= p7_add_8136_comb;
    p7_bit_slice_8137 <= p7_bit_slice_8137_comb;
    p7_ugt_8138 <= p7_ugt_8138_comb;
    p7_or_8139 <= p7_or_8139_comb;
    p7_ne_8141 <= p7_ne_8141_comb;
    p7_add_8142 <= p7_add_8142_comb;
    p7_bit_slice_8143 <= p7_bit_slice_8143_comb;
    p7_bd__1_sign <= p6_bd__1_sign;
    p7_result_sign__5 <= p6_result_sign__5;
    p7_result_sign__8 <= p6_result_sign__8;
    p7_result_sign__7 <= p6_result_sign__7;
    p7_eq_8148 <= p7_eq_8148_comb;
    p7_eq_8149 <= p7_eq_8149_comb;
    p7_eq_8150 <= p7_eq_8150_comb;
    p7_eq_8151 <= p7_eq_8151_comb;
    p7_ne_8156 <= p7_ne_8156_comb;
    p7_ne_8157 <= p7_ne_8157_comb;
    p7_ne_8158 <= p7_ne_8158_comb;
    p7_ne_8159 <= p7_ne_8159_comb;
    p7_in0_r_fraction__6 <= p6_in0_r_fraction__6;
    p7_in0_r_bexp__6 <= p6_in0_r_bexp__6;
    p7_in0_i_fraction__6 <= p6_in0_i_fraction__6;
    p7_in0_i_bexp__6 <= p6_in0_i_bexp__6;
    p7_in0_r_sign__2 <= p6_in0_r_sign__2;
    p7_in0_i_sign__2 <= p6_in0_i_sign__2;
  end

  // ===== Pipe stage 8:
  wire [27:0] p8_wide_x_comb;
  wire [7:0] p8_greater_exp_bexp_comb;
  wire [27:0] p8_wide_y_comb;
  wire [27:0] p8_wide_x__2_comb;
  wire [7:0] p8_greater_exp_bexp__1_comb;
  wire [27:0] p8_wide_y__2_comb;
  wire [7:0] p8_high_exp__32_comb;
  wire [7:0] p8_high_exp__33_comb;
  wire [7:0] p8_high_exp__34_comb;
  wire [7:0] p8_high_exp__35_comb;
  wire [27:0] p8_wide_x__1_comb;
  wire [7:0] p8_sub_8263_comb;
  wire [27:0] p8_wide_y__1_comb;
  wire [7:0] p8_sub_8265_comb;
  wire [27:0] p8_wide_x__3_comb;
  wire [7:0] p8_sub_8267_comb;
  wire [27:0] p8_wide_y__3_comb;
  wire [7:0] p8_sub_8269_comb;
  wire p8_eq_8300_comb;
  wire p8_eq_8301_comb;
  wire p8_eq_8302_comb;
  wire p8_eq_8303_comb;
  wire [27:0] p8_dropped_x_comb;
  wire [27:0] p8_dropped_y_comb;
  wire [27:0] p8_dropped_x__1_comb;
  wire [27:0] p8_dropped_y__1_comb;
  wire [7:0] p8_shift_x_comb;
  wire [7:0] p8_shift_y_comb;
  wire [7:0] p8_shift_x__1_comb;
  wire [7:0] p8_shift_y__1_comb;
  wire p8_sticky_x_comb;
  wire p8_sticky_y_comb;
  wire p8_sticky_x__1_comb;
  wire p8_sticky_y__1_comb;
  wire [27:0] p8_shifted_x_comb;
  wire [27:0] p8_shifted_y_comb;
  wire [27:0] p8_shifted_x__1_comb;
  wire [27:0] p8_shifted_y__1_comb;
  wire p8_greater_exp_sign_comb;
  wire p8_greater_exp_sign__1_comb;
  wire p8_and_8306_comb;
  wire p8_and_8307_comb;
  wire p8_and_8310_comb;
  wire p8_and_8311_comb;
  wire p8_has_pos_inf_comb;
  wire p8_has_pos_inf__1_comb;
  wire p8_and_8318_comb;
  wire p8_and_8319_comb;
  wire p8_and_8320_comb;
  wire p8_and_8321_comb;
  assign p8_wide_x_comb = {p7_or_8122, p7_literal_8123};
  assign p8_greater_exp_bexp_comb = p7_ugt_8127 ? p7_result_exp__8 : p7_result_exp__5;
  assign p8_wide_y_comb = {p7_or_8128, p7_literal_8129};
  assign p8_wide_x__2_comb = {p7_or_8133, p7_literal_8134};
  assign p8_greater_exp_bexp__1_comb = p7_ugt_8138 ? p7_result_exp__11 : p7_result_exp__12;
  assign p8_wide_y__2_comb = {p7_or_8139, p7_literal_8140};
  assign p8_high_exp__32_comb = 8'hff;
  assign p8_high_exp__33_comb = 8'hff;
  assign p8_high_exp__34_comb = 8'hff;
  assign p8_high_exp__35_comb = 8'hff;
  assign p8_wide_x__1_comb = p8_wide_x_comb & {28{p7_ne_8124}};
  assign p8_sub_8263_comb = {p7_add_8125, p7_bit_slice_8126} - p8_greater_exp_bexp_comb;
  assign p8_wide_y__1_comb = p8_wide_y_comb & {28{p7_ne_8130}};
  assign p8_sub_8265_comb = {p7_add_8131, p7_bit_slice_8132} - p8_greater_exp_bexp_comb;
  assign p8_wide_x__3_comb = p8_wide_x__2_comb & {28{p7_ne_8135}};
  assign p8_sub_8267_comb = {p7_add_8136, p7_bit_slice_8137} - p8_greater_exp_bexp__1_comb;
  assign p8_wide_y__3_comb = p8_wide_y__2_comb & {28{p7_ne_8141}};
  assign p8_sub_8269_comb = {p7_add_8142, p7_bit_slice_8143} - p8_greater_exp_bexp__1_comb;
  assign p8_eq_8300_comb = p7_result_exp__8 == p8_high_exp__32_comb;
  assign p8_eq_8301_comb = p7_result_exp__5 == p8_high_exp__33_comb;
  assign p8_eq_8302_comb = p7_result_exp__11 == p8_high_exp__34_comb;
  assign p8_eq_8303_comb = p7_result_exp__12 == p8_high_exp__35_comb;
  assign p8_dropped_x_comb = p8_sub_8263_comb >= 8'h1c ? 28'h000_0000 : p8_wide_x__1_comb << p8_sub_8263_comb;
  assign p8_dropped_y_comb = p8_sub_8265_comb >= 8'h1c ? 28'h000_0000 : p8_wide_y__1_comb << p8_sub_8265_comb;
  assign p8_dropped_x__1_comb = p8_sub_8267_comb >= 8'h1c ? 28'h000_0000 : p8_wide_x__3_comb << p8_sub_8267_comb;
  assign p8_dropped_y__1_comb = p8_sub_8269_comb >= 8'h1c ? 28'h000_0000 : p8_wide_y__3_comb << p8_sub_8269_comb;
  assign p8_shift_x_comb = p8_greater_exp_bexp_comb - p7_result_exp__8;
  assign p8_shift_y_comb = p8_greater_exp_bexp_comb - p7_result_exp__5;
  assign p8_shift_x__1_comb = p8_greater_exp_bexp__1_comb - p7_result_exp__11;
  assign p8_shift_y__1_comb = p8_greater_exp_bexp__1_comb - p7_result_exp__12;
  assign p8_sticky_x_comb = p8_dropped_x_comb[27:3] != 25'h000_0000;
  assign p8_sticky_y_comb = p8_dropped_y_comb[27:3] != 25'h000_0000;
  assign p8_sticky_x__1_comb = p8_dropped_x__1_comb[27:3] != 25'h000_0000;
  assign p8_sticky_y__1_comb = p8_dropped_y__1_comb[27:3] != 25'h000_0000;
  assign p8_shifted_x_comb = p8_shift_x_comb >= 8'h1c ? 28'h000_0000 : p8_wide_x__1_comb >> p8_shift_x_comb;
  assign p8_shifted_y_comb = p8_shift_y_comb >= 8'h1c ? 28'h000_0000 : p8_wide_y__1_comb >> p8_shift_y_comb;
  assign p8_shifted_x__1_comb = p8_shift_x__1_comb >= 8'h1c ? 28'h000_0000 : p8_wide_x__3_comb >> p8_shift_x__1_comb;
  assign p8_shifted_y__1_comb = p8_shift_y__1_comb >= 8'h1c ? 28'h000_0000 : p8_wide_y__3_comb >> p8_shift_y__1_comb;
  assign p8_greater_exp_sign_comb = p7_ugt_8127 ? p7_result_sign__5 : p7_bd__1_sign;
  assign p8_greater_exp_sign__1_comb = p7_ugt_8138 ? p7_result_sign__7 : p7_result_sign__8;
  assign p8_and_8306_comb = p8_eq_8300_comb & p7_eq_8148;
  assign p8_and_8307_comb = p8_eq_8301_comb & p7_eq_8149;
  assign p8_and_8310_comb = p8_eq_8302_comb & p7_eq_8150;
  assign p8_and_8311_comb = p8_eq_8303_comb & p7_eq_8151;
  assign p8_has_pos_inf_comb = ~(~(p8_eq_8300_comb & p7_eq_8148) | p7_result_sign__5) | ~(~(p8_eq_8301_comb & p7_eq_8149) | p7_bd__1_sign);
  assign p8_has_pos_inf__1_comb = ~(~(p8_eq_8302_comb & p7_eq_8150) | p7_result_sign__7) | ~(~(p8_eq_8303_comb & p7_eq_8151) | p7_result_sign__8);
  assign p8_and_8318_comb = p8_eq_8300_comb & p7_ne_8156;
  assign p8_and_8319_comb = p8_eq_8301_comb & p7_ne_8157;
  assign p8_and_8320_comb = p8_eq_8302_comb & p7_ne_8158;
  assign p8_and_8321_comb = p8_eq_8303_comb & p7_ne_8159;

  // Registers for pipe stage 8:
  reg [7:0] p8_greater_exp_bexp;
  reg [7:0] p8_greater_exp_bexp__1;
  reg p8_sticky_x;
  reg p8_sticky_y;
  reg p8_sticky_x__1;
  reg p8_sticky_y__1;
  reg p8_bd__1_sign;
  reg p8_result_sign__5;
  reg [27:0] p8_shifted_x;
  reg [27:0] p8_shifted_y;
  reg p8_result_sign__8;
  reg p8_result_sign__7;
  reg [27:0] p8_shifted_x__1;
  reg [27:0] p8_shifted_y__1;
  reg p8_greater_exp_sign;
  reg p8_greater_exp_sign__1;
  reg p8_and_8306;
  reg p8_and_8307;
  reg p8_and_8310;
  reg p8_and_8311;
  reg p8_has_pos_inf;
  reg p8_has_pos_inf__1;
  reg p8_and_8318;
  reg p8_and_8319;
  reg p8_and_8320;
  reg p8_and_8321;
  reg [22:0] p8_in0_r_fraction__6;
  reg [7:0] p8_in0_r_bexp__6;
  reg [22:0] p8_in0_i_fraction__6;
  reg [7:0] p8_in0_i_bexp__6;
  reg p8_in0_r_sign__2;
  reg p8_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p8_greater_exp_bexp <= p8_greater_exp_bexp_comb;
    p8_greater_exp_bexp__1 <= p8_greater_exp_bexp__1_comb;
    p8_sticky_x <= p8_sticky_x_comb;
    p8_sticky_y <= p8_sticky_y_comb;
    p8_sticky_x__1 <= p8_sticky_x__1_comb;
    p8_sticky_y__1 <= p8_sticky_y__1_comb;
    p8_bd__1_sign <= p7_bd__1_sign;
    p8_result_sign__5 <= p7_result_sign__5;
    p8_shifted_x <= p8_shifted_x_comb;
    p8_shifted_y <= p8_shifted_y_comb;
    p8_result_sign__8 <= p7_result_sign__8;
    p8_result_sign__7 <= p7_result_sign__7;
    p8_shifted_x__1 <= p8_shifted_x__1_comb;
    p8_shifted_y__1 <= p8_shifted_y__1_comb;
    p8_greater_exp_sign <= p8_greater_exp_sign_comb;
    p8_greater_exp_sign__1 <= p8_greater_exp_sign__1_comb;
    p8_and_8306 <= p8_and_8306_comb;
    p8_and_8307 <= p8_and_8307_comb;
    p8_and_8310 <= p8_and_8310_comb;
    p8_and_8311 <= p8_and_8311_comb;
    p8_has_pos_inf <= p8_has_pos_inf_comb;
    p8_has_pos_inf__1 <= p8_has_pos_inf__1_comb;
    p8_and_8318 <= p8_and_8318_comb;
    p8_and_8319 <= p8_and_8319_comb;
    p8_and_8320 <= p8_and_8320_comb;
    p8_and_8321 <= p8_and_8321_comb;
    p8_in0_r_fraction__6 <= p7_in0_r_fraction__6;
    p8_in0_r_bexp__6 <= p7_in0_r_bexp__6;
    p8_in0_i_fraction__6 <= p7_in0_i_fraction__6;
    p8_in0_i_bexp__6 <= p7_in0_i_bexp__6;
    p8_in0_r_sign__2 <= p7_in0_r_sign__2;
    p8_in0_i_sign__2 <= p7_in0_i_sign__2;
  end

  // ===== Pipe stage 9:
  wire [27:0] p9_addend_x_comb;
  wire [27:0] p9_addend_y_comb;
  wire [27:0] p9_addend_x__2_comb;
  wire [27:0] p9_addend_y__2_comb;
  wire p9_has_neg_inf_comb;
  wire p9_has_neg_inf__1_comb;
  wire [27:0] p9_addend_x__1_comb;
  wire [27:0] p9_addend_y__1_comb;
  wire [27:0] p9_addend_x__3_comb;
  wire [27:0] p9_addend_y__3_comb;
  wire p9_nor_8416_comb;
  wire p9_nor_8418_comb;
  wire p9_is_result_nan__5_comb;
  wire p9_is_operand_inf_comb;
  wire p9_is_result_nan__6_comb;
  wire p9_is_operand_inf__1_comb;
  wire p9_not_8424_comb;
  wire p9_not_8425_comb;
  assign p9_addend_x_comb = p8_shifted_x | {27'h000_0000, p8_sticky_x};
  assign p9_addend_y_comb = p8_shifted_y | {27'h000_0000, p8_sticky_y};
  assign p9_addend_x__2_comb = p8_shifted_x__1 | {27'h000_0000, p8_sticky_x__1};
  assign p9_addend_y__2_comb = p8_shifted_y__1 | {27'h000_0000, p8_sticky_y__1};
  assign p9_has_neg_inf_comb = p8_and_8306 & p8_result_sign__5 | p8_and_8307 & p8_bd__1_sign;
  assign p9_has_neg_inf__1_comb = p8_and_8310 & p8_result_sign__7 | p8_and_8311 & p8_result_sign__8;
  assign p9_addend_x__1_comb = p8_result_sign__5 ^ p8_greater_exp_sign ? -p9_addend_x_comb : p9_addend_x_comb;
  assign p9_addend_y__1_comb = p8_bd__1_sign ^ p8_greater_exp_sign ? -p9_addend_y_comb : p9_addend_y_comb;
  assign p9_addend_x__3_comb = p8_result_sign__7 ^ p8_greater_exp_sign__1 ? -p9_addend_x__2_comb : p9_addend_x__2_comb;
  assign p9_addend_y__3_comb = p8_result_sign__8 ^ p8_greater_exp_sign__1 ? -p9_addend_y__2_comb : p9_addend_y__2_comb;
  assign p9_nor_8416_comb = ~(p8_and_8306 | p8_and_8307);
  assign p9_nor_8418_comb = ~(p8_and_8310 | p8_and_8311);
  assign p9_is_result_nan__5_comb = p8_and_8318 | p8_and_8319 | p8_has_pos_inf & p9_has_neg_inf_comb;
  assign p9_is_operand_inf_comb = p8_and_8306 | p8_and_8307;
  assign p9_is_result_nan__6_comb = p8_and_8320 | p8_and_8321 | p8_has_pos_inf__1 & p9_has_neg_inf__1_comb;
  assign p9_is_operand_inf__1_comb = p8_and_8310 | p8_and_8311;
  assign p9_not_8424_comb = ~p8_has_pos_inf;
  assign p9_not_8425_comb = ~p8_has_pos_inf__1;

  // Registers for pipe stage 9:
  reg [7:0] p9_greater_exp_bexp;
  reg [7:0] p9_greater_exp_bexp__1;
  reg p9_greater_exp_sign;
  reg p9_greater_exp_sign__1;
  reg [27:0] p9_addend_x__1;
  reg [27:0] p9_addend_y__1;
  reg [27:0] p9_addend_x__3;
  reg [27:0] p9_addend_y__3;
  reg p9_nor_8416;
  reg p9_nor_8418;
  reg p9_is_result_nan__5;
  reg p9_is_operand_inf;
  reg p9_is_result_nan__6;
  reg p9_is_operand_inf__1;
  reg [22:0] p9_in0_r_fraction__6;
  reg [7:0] p9_in0_r_bexp__6;
  reg [22:0] p9_in0_i_fraction__6;
  reg [7:0] p9_in0_i_bexp__6;
  reg p9_not_8424;
  reg p9_not_8425;
  reg p9_in0_r_sign__2;
  reg p9_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p9_greater_exp_bexp <= p8_greater_exp_bexp;
    p9_greater_exp_bexp__1 <= p8_greater_exp_bexp__1;
    p9_greater_exp_sign <= p8_greater_exp_sign;
    p9_greater_exp_sign__1 <= p8_greater_exp_sign__1;
    p9_addend_x__1 <= p9_addend_x__1_comb;
    p9_addend_y__1 <= p9_addend_y__1_comb;
    p9_addend_x__3 <= p9_addend_x__3_comb;
    p9_addend_y__3 <= p9_addend_y__3_comb;
    p9_nor_8416 <= p9_nor_8416_comb;
    p9_nor_8418 <= p9_nor_8418_comb;
    p9_is_result_nan__5 <= p9_is_result_nan__5_comb;
    p9_is_operand_inf <= p9_is_operand_inf_comb;
    p9_is_result_nan__6 <= p9_is_result_nan__6_comb;
    p9_is_operand_inf__1 <= p9_is_operand_inf__1_comb;
    p9_in0_r_fraction__6 <= p8_in0_r_fraction__6;
    p9_in0_r_bexp__6 <= p8_in0_r_bexp__6;
    p9_in0_i_fraction__6 <= p8_in0_i_fraction__6;
    p9_in0_i_bexp__6 <= p8_in0_i_bexp__6;
    p9_not_8424 <= p9_not_8424_comb;
    p9_not_8425 <= p9_not_8425_comb;
    p9_in0_r_sign__2 <= p8_in0_r_sign__2;
    p9_in0_i_sign__2 <= p8_in0_i_sign__2;
  end

  // ===== Pipe stage 10:
  wire [28:0] p10_fraction__33_comb;
  wire [28:0] p10_fraction__34_comb;
  wire p10_fraction_is_zero_comb;
  wire p10_fraction_is_zero__1_comb;
  wire [27:0] p10_abs_fraction_comb;
  wire [27:0] p10_abs_fraction__1_comb;
  wire p10_ne_8486_comb;
  wire p10_ne_8487_comb;
  wire p10_nor_8496_comb;
  wire p10_nor_8497_comb;
  wire p10_nor_8498_comb;
  wire p10_nor_8499_comb;
  assign p10_fraction__33_comb = {{1{p9_addend_x__1[27]}}, p9_addend_x__1} + {{1{p9_addend_y__1[27]}}, p9_addend_y__1};
  assign p10_fraction__34_comb = {{1{p9_addend_x__3[27]}}, p9_addend_x__3} + {{1{p9_addend_y__3[27]}}, p9_addend_y__3};
  assign p10_fraction_is_zero_comb = p10_fraction__33_comb == 29'h0000_0000;
  assign p10_fraction_is_zero__1_comb = p10_fraction__34_comb == 29'h0000_0000;
  assign p10_abs_fraction_comb = p10_fraction__33_comb[28] ? -p10_fraction__33_comb[27:0] : p10_fraction__33_comb[27:0];
  assign p10_abs_fraction__1_comb = p10_fraction__34_comb[28] ? -p10_fraction__34_comb[27:0] : p10_fraction__34_comb[27:0];
  assign p10_ne_8486_comb = p10_fraction__33_comb != 29'h0000_0000;
  assign p10_ne_8487_comb = p10_fraction__34_comb != 29'h0000_0000;
  assign p10_nor_8496_comb = ~(~p10_fraction__33_comb[28] | p9_greater_exp_sign);
  assign p10_nor_8497_comb = ~(p10_fraction__33_comb[28] | p10_fraction_is_zero_comb | ~p9_greater_exp_sign);
  assign p10_nor_8498_comb = ~(~p10_fraction__34_comb[28] | p9_greater_exp_sign__1);
  assign p10_nor_8499_comb = ~(p10_fraction__34_comb[28] | p10_fraction_is_zero__1_comb | ~p9_greater_exp_sign__1);

  // Registers for pipe stage 10:
  reg [7:0] p10_greater_exp_bexp;
  reg [7:0] p10_greater_exp_bexp__1;
  reg [27:0] p10_abs_fraction;
  reg [27:0] p10_abs_fraction__1;
  reg p10_ne_8486;
  reg p10_ne_8487;
  reg p10_nor_8416;
  reg p10_nor_8418;
  reg p10_is_result_nan__5;
  reg p10_is_operand_inf;
  reg p10_is_result_nan__6;
  reg p10_is_operand_inf__1;
  reg [22:0] p10_in0_r_fraction__6;
  reg [7:0] p10_in0_r_bexp__6;
  reg [22:0] p10_in0_i_fraction__6;
  reg [7:0] p10_in0_i_bexp__6;
  reg p10_nor_8496;
  reg p10_nor_8497;
  reg p10_nor_8498;
  reg p10_nor_8499;
  reg p10_not_8424;
  reg p10_not_8425;
  reg p10_in0_r_sign__2;
  reg p10_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p10_greater_exp_bexp <= p9_greater_exp_bexp;
    p10_greater_exp_bexp__1 <= p9_greater_exp_bexp__1;
    p10_abs_fraction <= p10_abs_fraction_comb;
    p10_abs_fraction__1 <= p10_abs_fraction__1_comb;
    p10_ne_8486 <= p10_ne_8486_comb;
    p10_ne_8487 <= p10_ne_8487_comb;
    p10_nor_8416 <= p9_nor_8416;
    p10_nor_8418 <= p9_nor_8418;
    p10_is_result_nan__5 <= p9_is_result_nan__5;
    p10_is_operand_inf <= p9_is_operand_inf;
    p10_is_result_nan__6 <= p9_is_result_nan__6;
    p10_is_operand_inf__1 <= p9_is_operand_inf__1;
    p10_in0_r_fraction__6 <= p9_in0_r_fraction__6;
    p10_in0_r_bexp__6 <= p9_in0_r_bexp__6;
    p10_in0_i_fraction__6 <= p9_in0_i_fraction__6;
    p10_in0_i_bexp__6 <= p9_in0_i_bexp__6;
    p10_nor_8496 <= p10_nor_8496_comb;
    p10_nor_8497 <= p10_nor_8497_comb;
    p10_nor_8498 <= p10_nor_8498_comb;
    p10_nor_8499 <= p10_nor_8499_comb;
    p10_not_8424 <= p9_not_8424;
    p10_not_8425 <= p9_not_8425;
    p10_in0_r_sign__2 <= p9_in0_r_sign__2;
    p10_in0_i_sign__2 <= p9_in0_i_sign__2;
  end

  // ===== Pipe stage 11:
  wire [27:0] p11_reverse_8548_comb;
  wire [27:0] p11_reverse_8549_comb;
  wire [28:0] p11_one_hot_8550_comb;
  wire [28:0] p11_one_hot_8551_comb;
  wire [4:0] p11_encode_8552_comb;
  wire [4:0] p11_encode_8553_comb;
  wire p11_result_sign__9_comb;
  wire p11_result_sign__11_comb;
  wire p11_result_sign__10_comb;
  wire p11_result_sign__12_comb;
  wire p11_cancel_comb;
  wire p11_cancel__1_comb;
  wire p11_result_sign__13_comb;
  wire p11_result_sign__14_comb;
  assign p11_reverse_8548_comb = {p10_abs_fraction[0], p10_abs_fraction[1], p10_abs_fraction[2], p10_abs_fraction[3], p10_abs_fraction[4], p10_abs_fraction[5], p10_abs_fraction[6], p10_abs_fraction[7], p10_abs_fraction[8], p10_abs_fraction[9], p10_abs_fraction[10], p10_abs_fraction[11], p10_abs_fraction[12], p10_abs_fraction[13], p10_abs_fraction[14], p10_abs_fraction[15], p10_abs_fraction[16], p10_abs_fraction[17], p10_abs_fraction[18], p10_abs_fraction[19], p10_abs_fraction[20], p10_abs_fraction[21], p10_abs_fraction[22], p10_abs_fraction[23], p10_abs_fraction[24], p10_abs_fraction[25], p10_abs_fraction[26], p10_abs_fraction[27]};
  assign p11_reverse_8549_comb = {p10_abs_fraction__1[0], p10_abs_fraction__1[1], p10_abs_fraction__1[2], p10_abs_fraction__1[3], p10_abs_fraction__1[4], p10_abs_fraction__1[5], p10_abs_fraction__1[6], p10_abs_fraction__1[7], p10_abs_fraction__1[8], p10_abs_fraction__1[9], p10_abs_fraction__1[10], p10_abs_fraction__1[11], p10_abs_fraction__1[12], p10_abs_fraction__1[13], p10_abs_fraction__1[14], p10_abs_fraction__1[15], p10_abs_fraction__1[16], p10_abs_fraction__1[17], p10_abs_fraction__1[18], p10_abs_fraction__1[19], p10_abs_fraction__1[20], p10_abs_fraction__1[21], p10_abs_fraction__1[22], p10_abs_fraction__1[23], p10_abs_fraction__1[24], p10_abs_fraction__1[25], p10_abs_fraction__1[26], p10_abs_fraction__1[27]};
  assign p11_one_hot_8550_comb = {p11_reverse_8548_comb[27:0] == 28'h000_0000, p11_reverse_8548_comb[27] && p11_reverse_8548_comb[26:0] == 27'h000_0000, p11_reverse_8548_comb[26] && p11_reverse_8548_comb[25:0] == 26'h000_0000, p11_reverse_8548_comb[25] && p11_reverse_8548_comb[24:0] == 25'h000_0000, p11_reverse_8548_comb[24] && p11_reverse_8548_comb[23:0] == 24'h00_0000, p11_reverse_8548_comb[23] && p11_reverse_8548_comb[22:0] == 23'h00_0000, p11_reverse_8548_comb[22] && p11_reverse_8548_comb[21:0] == 22'h00_0000, p11_reverse_8548_comb[21] && p11_reverse_8548_comb[20:0] == 21'h00_0000, p11_reverse_8548_comb[20] && p11_reverse_8548_comb[19:0] == 20'h0_0000, p11_reverse_8548_comb[19] && p11_reverse_8548_comb[18:0] == 19'h0_0000, p11_reverse_8548_comb[18] && p11_reverse_8548_comb[17:0] == 18'h0_0000, p11_reverse_8548_comb[17] && p11_reverse_8548_comb[16:0] == 17'h0_0000, p11_reverse_8548_comb[16] && p11_reverse_8548_comb[15:0] == 16'h0000, p11_reverse_8548_comb[15] && p11_reverse_8548_comb[14:0] == 15'h0000, p11_reverse_8548_comb[14] && p11_reverse_8548_comb[13:0] == 14'h0000, p11_reverse_8548_comb[13] && p11_reverse_8548_comb[12:0] == 13'h0000, p11_reverse_8548_comb[12] && p11_reverse_8548_comb[11:0] == 12'h000, p11_reverse_8548_comb[11] && p11_reverse_8548_comb[10:0] == 11'h000, p11_reverse_8548_comb[10] && p11_reverse_8548_comb[9:0] == 10'h000, p11_reverse_8548_comb[9] && p11_reverse_8548_comb[8:0] == 9'h000, p11_reverse_8548_comb[8] && p11_reverse_8548_comb[7:0] == 8'h00, p11_reverse_8548_comb[7] && p11_reverse_8548_comb[6:0] == 7'h00, p11_reverse_8548_comb[6] && p11_reverse_8548_comb[5:0] == 6'h00, p11_reverse_8548_comb[5] && p11_reverse_8548_comb[4:0] == 5'h00, p11_reverse_8548_comb[4] && p11_reverse_8548_comb[3:0] == 4'h0, p11_reverse_8548_comb[3] && p11_reverse_8548_comb[2:0] == 3'h0, p11_reverse_8548_comb[2] && p11_reverse_8548_comb[1:0] == 2'h0, p11_reverse_8548_comb[1] && !p11_reverse_8548_comb[0], p11_reverse_8548_comb[0]};
  assign p11_one_hot_8551_comb = {p11_reverse_8549_comb[27:0] == 28'h000_0000, p11_reverse_8549_comb[27] && p11_reverse_8549_comb[26:0] == 27'h000_0000, p11_reverse_8549_comb[26] && p11_reverse_8549_comb[25:0] == 26'h000_0000, p11_reverse_8549_comb[25] && p11_reverse_8549_comb[24:0] == 25'h000_0000, p11_reverse_8549_comb[24] && p11_reverse_8549_comb[23:0] == 24'h00_0000, p11_reverse_8549_comb[23] && p11_reverse_8549_comb[22:0] == 23'h00_0000, p11_reverse_8549_comb[22] && p11_reverse_8549_comb[21:0] == 22'h00_0000, p11_reverse_8549_comb[21] && p11_reverse_8549_comb[20:0] == 21'h00_0000, p11_reverse_8549_comb[20] && p11_reverse_8549_comb[19:0] == 20'h0_0000, p11_reverse_8549_comb[19] && p11_reverse_8549_comb[18:0] == 19'h0_0000, p11_reverse_8549_comb[18] && p11_reverse_8549_comb[17:0] == 18'h0_0000, p11_reverse_8549_comb[17] && p11_reverse_8549_comb[16:0] == 17'h0_0000, p11_reverse_8549_comb[16] && p11_reverse_8549_comb[15:0] == 16'h0000, p11_reverse_8549_comb[15] && p11_reverse_8549_comb[14:0] == 15'h0000, p11_reverse_8549_comb[14] && p11_reverse_8549_comb[13:0] == 14'h0000, p11_reverse_8549_comb[13] && p11_reverse_8549_comb[12:0] == 13'h0000, p11_reverse_8549_comb[12] && p11_reverse_8549_comb[11:0] == 12'h000, p11_reverse_8549_comb[11] && p11_reverse_8549_comb[10:0] == 11'h000, p11_reverse_8549_comb[10] && p11_reverse_8549_comb[9:0] == 10'h000, p11_reverse_8549_comb[9] && p11_reverse_8549_comb[8:0] == 9'h000, p11_reverse_8549_comb[8] && p11_reverse_8549_comb[7:0] == 8'h00, p11_reverse_8549_comb[7] && p11_reverse_8549_comb[6:0] == 7'h00, p11_reverse_8549_comb[6] && p11_reverse_8549_comb[5:0] == 6'h00, p11_reverse_8549_comb[5] && p11_reverse_8549_comb[4:0] == 5'h00, p11_reverse_8549_comb[4] && p11_reverse_8549_comb[3:0] == 4'h0, p11_reverse_8549_comb[3] && p11_reverse_8549_comb[2:0] == 3'h0, p11_reverse_8549_comb[2] && p11_reverse_8549_comb[1:0] == 2'h0, p11_reverse_8549_comb[1] && !p11_reverse_8549_comb[0], p11_reverse_8549_comb[0]};
  assign p11_encode_8552_comb = {p11_one_hot_8550_comb[16] | p11_one_hot_8550_comb[17] | p11_one_hot_8550_comb[18] | p11_one_hot_8550_comb[19] | p11_one_hot_8550_comb[20] | p11_one_hot_8550_comb[21] | p11_one_hot_8550_comb[22] | p11_one_hot_8550_comb[23] | p11_one_hot_8550_comb[24] | p11_one_hot_8550_comb[25] | p11_one_hot_8550_comb[26] | p11_one_hot_8550_comb[27] | p11_one_hot_8550_comb[28], p11_one_hot_8550_comb[8] | p11_one_hot_8550_comb[9] | p11_one_hot_8550_comb[10] | p11_one_hot_8550_comb[11] | p11_one_hot_8550_comb[12] | p11_one_hot_8550_comb[13] | p11_one_hot_8550_comb[14] | p11_one_hot_8550_comb[15] | p11_one_hot_8550_comb[24] | p11_one_hot_8550_comb[25] | p11_one_hot_8550_comb[26] | p11_one_hot_8550_comb[27] | p11_one_hot_8550_comb[28], p11_one_hot_8550_comb[4] | p11_one_hot_8550_comb[5] | p11_one_hot_8550_comb[6] | p11_one_hot_8550_comb[7] | p11_one_hot_8550_comb[12] | p11_one_hot_8550_comb[13] | p11_one_hot_8550_comb[14] | p11_one_hot_8550_comb[15] | p11_one_hot_8550_comb[20] | p11_one_hot_8550_comb[21] | p11_one_hot_8550_comb[22] | p11_one_hot_8550_comb[23] | p11_one_hot_8550_comb[28], p11_one_hot_8550_comb[2] | p11_one_hot_8550_comb[3] | p11_one_hot_8550_comb[6] | p11_one_hot_8550_comb[7] | p11_one_hot_8550_comb[10] | p11_one_hot_8550_comb[11] | p11_one_hot_8550_comb[14] | p11_one_hot_8550_comb[15] | p11_one_hot_8550_comb[18] | p11_one_hot_8550_comb[19] | p11_one_hot_8550_comb[22] | p11_one_hot_8550_comb[23] | p11_one_hot_8550_comb[26] | p11_one_hot_8550_comb[27], p11_one_hot_8550_comb[1] | p11_one_hot_8550_comb[3] | p11_one_hot_8550_comb[5] | p11_one_hot_8550_comb[7] | p11_one_hot_8550_comb[9] | p11_one_hot_8550_comb[11] | p11_one_hot_8550_comb[13] | p11_one_hot_8550_comb[15] | p11_one_hot_8550_comb[17] | p11_one_hot_8550_comb[19] | p11_one_hot_8550_comb[21] | p11_one_hot_8550_comb[23] | p11_one_hot_8550_comb[25] | p11_one_hot_8550_comb[27]};
  assign p11_encode_8553_comb = {p11_one_hot_8551_comb[16] | p11_one_hot_8551_comb[17] | p11_one_hot_8551_comb[18] | p11_one_hot_8551_comb[19] | p11_one_hot_8551_comb[20] | p11_one_hot_8551_comb[21] | p11_one_hot_8551_comb[22] | p11_one_hot_8551_comb[23] | p11_one_hot_8551_comb[24] | p11_one_hot_8551_comb[25] | p11_one_hot_8551_comb[26] | p11_one_hot_8551_comb[27] | p11_one_hot_8551_comb[28], p11_one_hot_8551_comb[8] | p11_one_hot_8551_comb[9] | p11_one_hot_8551_comb[10] | p11_one_hot_8551_comb[11] | p11_one_hot_8551_comb[12] | p11_one_hot_8551_comb[13] | p11_one_hot_8551_comb[14] | p11_one_hot_8551_comb[15] | p11_one_hot_8551_comb[24] | p11_one_hot_8551_comb[25] | p11_one_hot_8551_comb[26] | p11_one_hot_8551_comb[27] | p11_one_hot_8551_comb[28], p11_one_hot_8551_comb[4] | p11_one_hot_8551_comb[5] | p11_one_hot_8551_comb[6] | p11_one_hot_8551_comb[7] | p11_one_hot_8551_comb[12] | p11_one_hot_8551_comb[13] | p11_one_hot_8551_comb[14] | p11_one_hot_8551_comb[15] | p11_one_hot_8551_comb[20] | p11_one_hot_8551_comb[21] | p11_one_hot_8551_comb[22] | p11_one_hot_8551_comb[23] | p11_one_hot_8551_comb[28], p11_one_hot_8551_comb[2] | p11_one_hot_8551_comb[3] | p11_one_hot_8551_comb[6] | p11_one_hot_8551_comb[7] | p11_one_hot_8551_comb[10] | p11_one_hot_8551_comb[11] | p11_one_hot_8551_comb[14] | p11_one_hot_8551_comb[15] | p11_one_hot_8551_comb[18] | p11_one_hot_8551_comb[19] | p11_one_hot_8551_comb[22] | p11_one_hot_8551_comb[23] | p11_one_hot_8551_comb[26] | p11_one_hot_8551_comb[27], p11_one_hot_8551_comb[1] | p11_one_hot_8551_comb[3] | p11_one_hot_8551_comb[5] | p11_one_hot_8551_comb[7] | p11_one_hot_8551_comb[9] | p11_one_hot_8551_comb[11] | p11_one_hot_8551_comb[13] | p11_one_hot_8551_comb[15] | p11_one_hot_8551_comb[17] | p11_one_hot_8551_comb[19] | p11_one_hot_8551_comb[21] | p11_one_hot_8551_comb[23] | p11_one_hot_8551_comb[25] | p11_one_hot_8551_comb[27]};
  assign p11_result_sign__9_comb = p10_nor_8496 | p10_nor_8497;
  assign p11_result_sign__11_comb = p10_nor_8498 | p10_nor_8499;
  assign p11_result_sign__10_comb = p10_is_operand_inf ? p10_not_8424 : p11_result_sign__9_comb;
  assign p11_result_sign__12_comb = p10_is_operand_inf__1 ? p10_not_8425 : p11_result_sign__11_comb;
  assign p11_cancel_comb = p11_encode_8552_comb[1] | p11_encode_8552_comb[2] | p11_encode_8552_comb[3] | p11_encode_8552_comb[4];
  assign p11_cancel__1_comb = p11_encode_8553_comb[1] | p11_encode_8553_comb[2] | p11_encode_8553_comb[3] | p11_encode_8553_comb[4];
  assign p11_result_sign__13_comb = ~p10_is_result_nan__5 & p11_result_sign__10_comb;
  assign p11_result_sign__14_comb = ~p10_is_result_nan__6 & p11_result_sign__12_comb;

  // Registers for pipe stage 11:
  reg [7:0] p11_greater_exp_bexp;
  reg [7:0] p11_greater_exp_bexp__1;
  reg [27:0] p11_abs_fraction;
  reg [27:0] p11_abs_fraction__1;
  reg [4:0] p11_encode_8552;
  reg [4:0] p11_encode_8553;
  reg p11_cancel;
  reg p11_cancel__1;
  reg p11_ne_8486;
  reg p11_ne_8487;
  reg p11_nor_8416;
  reg p11_nor_8418;
  reg p11_is_result_nan__5;
  reg p11_is_operand_inf;
  reg p11_is_result_nan__6;
  reg p11_is_operand_inf__1;
  reg [22:0] p11_in0_r_fraction__6;
  reg [7:0] p11_in0_r_bexp__6;
  reg [22:0] p11_in0_i_fraction__6;
  reg [7:0] p11_in0_i_bexp__6;
  reg p11_result_sign__13;
  reg p11_result_sign__14;
  reg p11_in0_r_sign__2;
  reg p11_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p11_greater_exp_bexp <= p10_greater_exp_bexp;
    p11_greater_exp_bexp__1 <= p10_greater_exp_bexp__1;
    p11_abs_fraction <= p10_abs_fraction;
    p11_abs_fraction__1 <= p10_abs_fraction__1;
    p11_encode_8552 <= p11_encode_8552_comb;
    p11_encode_8553 <= p11_encode_8553_comb;
    p11_cancel <= p11_cancel_comb;
    p11_cancel__1 <= p11_cancel__1_comb;
    p11_ne_8486 <= p10_ne_8486;
    p11_ne_8487 <= p10_ne_8487;
    p11_nor_8416 <= p10_nor_8416;
    p11_nor_8418 <= p10_nor_8418;
    p11_is_result_nan__5 <= p10_is_result_nan__5;
    p11_is_operand_inf <= p10_is_operand_inf;
    p11_is_result_nan__6 <= p10_is_result_nan__6;
    p11_is_operand_inf__1 <= p10_is_operand_inf__1;
    p11_in0_r_fraction__6 <= p10_in0_r_fraction__6;
    p11_in0_r_bexp__6 <= p10_in0_r_bexp__6;
    p11_in0_i_fraction__6 <= p10_in0_i_fraction__6;
    p11_in0_i_bexp__6 <= p10_in0_i_bexp__6;
    p11_result_sign__13 <= p11_result_sign__13_comb;
    p11_result_sign__14 <= p11_result_sign__14_comb;
    p11_in0_r_sign__2 <= p10_in0_r_sign__2;
    p11_in0_i_sign__2 <= p10_in0_i_sign__2;
  end

  // ===== Pipe stage 12:
  wire p12_carry_bit_comb;
  wire p12_carry_bit__1_comb;
  wire [27:0] p12_leading_zeroes_comb;
  wire [27:0] p12_leading_zeroes__1_comb;
  wire [26:0] p12_carry_fraction_comb;
  wire [27:0] p12_add_8642_comb;
  wire [26:0] p12_carry_fraction__2_comb;
  wire [27:0] p12_add_8649_comb;
  wire [2:0] p12_concat_8650_comb;
  wire [26:0] p12_carry_fraction__1_comb;
  wire [26:0] p12_cancel_fraction_comb;
  wire [2:0] p12_concat_8653_comb;
  wire [26:0] p12_carry_fraction__3_comb;
  wire [26:0] p12_cancel_fraction__1_comb;
  wire [26:0] p12_shifted_fraction_comb;
  wire [26:0] p12_shifted_fraction__1_comb;
  assign p12_carry_bit_comb = p11_abs_fraction[27];
  assign p12_carry_bit__1_comb = p11_abs_fraction__1[27];
  assign p12_leading_zeroes_comb = {23'h00_0000, p11_encode_8552};
  assign p12_leading_zeroes__1_comb = {23'h00_0000, p11_encode_8553};
  assign p12_carry_fraction_comb = p11_abs_fraction[27:1];
  assign p12_add_8642_comb = p12_leading_zeroes_comb + 28'hfff_ffff;
  assign p12_carry_fraction__2_comb = p11_abs_fraction__1[27:1];
  assign p12_add_8649_comb = p12_leading_zeroes__1_comb + 28'hfff_ffff;
  assign p12_concat_8650_comb = {~p12_carry_bit_comb & ~p11_cancel, ~p12_carry_bit_comb & p11_cancel, p12_carry_bit_comb & ~p11_cancel};
  assign p12_carry_fraction__1_comb = p12_carry_fraction_comb | {26'h000_0000, p11_abs_fraction[0]};
  assign p12_cancel_fraction_comb = p12_add_8642_comb >= 28'h000_001b ? 27'h000_0000 : p11_abs_fraction[26:0] << p12_add_8642_comb;
  assign p12_concat_8653_comb = {~p12_carry_bit__1_comb & ~p11_cancel__1, ~p12_carry_bit__1_comb & p11_cancel__1, p12_carry_bit__1_comb & ~p11_cancel__1};
  assign p12_carry_fraction__3_comb = p12_carry_fraction__2_comb | {26'h000_0000, p11_abs_fraction__1[0]};
  assign p12_cancel_fraction__1_comb = p12_add_8649_comb >= 28'h000_001b ? 27'h000_0000 : p11_abs_fraction__1[26:0] << p12_add_8649_comb;
  assign p12_shifted_fraction_comb = p12_carry_fraction__1_comb & {27{p12_concat_8650_comb[0]}} | p12_cancel_fraction_comb & {27{p12_concat_8650_comb[1]}} | p11_abs_fraction[26:0] & {27{p12_concat_8650_comb[2]}};
  assign p12_shifted_fraction__1_comb = p12_carry_fraction__3_comb & {27{p12_concat_8653_comb[0]}} | p12_cancel_fraction__1_comb & {27{p12_concat_8653_comb[1]}} | p11_abs_fraction__1[26:0] & {27{p12_concat_8653_comb[2]}};

  // Registers for pipe stage 12:
  reg [7:0] p12_greater_exp_bexp;
  reg [7:0] p12_greater_exp_bexp__1;
  reg [4:0] p12_encode_8552;
  reg [4:0] p12_encode_8553;
  reg [26:0] p12_shifted_fraction;
  reg [26:0] p12_shifted_fraction__1;
  reg p12_ne_8486;
  reg p12_ne_8487;
  reg p12_nor_8416;
  reg p12_nor_8418;
  reg p12_is_result_nan__5;
  reg p12_is_operand_inf;
  reg p12_is_result_nan__6;
  reg p12_is_operand_inf__1;
  reg [22:0] p12_in0_r_fraction__6;
  reg [7:0] p12_in0_r_bexp__6;
  reg [22:0] p12_in0_i_fraction__6;
  reg [7:0] p12_in0_i_bexp__6;
  reg p12_result_sign__13;
  reg p12_result_sign__14;
  reg p12_in0_r_sign__2;
  reg p12_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p12_greater_exp_bexp <= p11_greater_exp_bexp;
    p12_greater_exp_bexp__1 <= p11_greater_exp_bexp__1;
    p12_encode_8552 <= p11_encode_8552;
    p12_encode_8553 <= p11_encode_8553;
    p12_shifted_fraction <= p12_shifted_fraction_comb;
    p12_shifted_fraction__1 <= p12_shifted_fraction__1_comb;
    p12_ne_8486 <= p11_ne_8486;
    p12_ne_8487 <= p11_ne_8487;
    p12_nor_8416 <= p11_nor_8416;
    p12_nor_8418 <= p11_nor_8418;
    p12_is_result_nan__5 <= p11_is_result_nan__5;
    p12_is_operand_inf <= p11_is_operand_inf;
    p12_is_result_nan__6 <= p11_is_result_nan__6;
    p12_is_operand_inf__1 <= p11_is_operand_inf__1;
    p12_in0_r_fraction__6 <= p11_in0_r_fraction__6;
    p12_in0_r_bexp__6 <= p11_in0_r_bexp__6;
    p12_in0_i_fraction__6 <= p11_in0_i_fraction__6;
    p12_in0_i_bexp__6 <= p11_in0_i_bexp__6;
    p12_result_sign__13 <= p11_result_sign__13;
    p12_result_sign__14 <= p11_result_sign__14;
    p12_in0_r_sign__2 <= p11_in0_r_sign__2;
    p12_in0_i_sign__2 <= p11_in0_i_sign__2;
  end

  // ===== Pipe stage 13:
  wire [2:0] p13_normal_chunk_comb;
  wire [1:0] p13_half_way_chunk_comb;
  wire [2:0] p13_normal_chunk__1_comb;
  wire [1:0] p13_half_way_chunk__1_comb;
  wire [24:0] p13_add_8721_comb;
  wire [24:0] p13_add_8725_comb;
  wire p13_do_round_up__5_comb;
  wire p13_do_round_up__6_comb;
  wire [27:0] p13_rounded_fraction_comb;
  wire [27:0] p13_rounded_fraction__1_comb;
  assign p13_normal_chunk_comb = p12_shifted_fraction[2:0];
  assign p13_half_way_chunk_comb = p12_shifted_fraction[3:2];
  assign p13_normal_chunk__1_comb = p12_shifted_fraction__1[2:0];
  assign p13_half_way_chunk__1_comb = p12_shifted_fraction__1[3:2];
  assign p13_add_8721_comb = {1'h0, p12_shifted_fraction[26:3]} + 25'h000_0001;
  assign p13_add_8725_comb = {1'h0, p12_shifted_fraction__1[26:3]} + 25'h000_0001;
  assign p13_do_round_up__5_comb = p13_normal_chunk_comb > 3'h4 | p13_half_way_chunk_comb == 2'h3;
  assign p13_do_round_up__6_comb = p13_normal_chunk__1_comb > 3'h4 | p13_half_way_chunk__1_comb == 2'h3;
  assign p13_rounded_fraction_comb = p13_do_round_up__5_comb ? {p13_add_8721_comb, p13_normal_chunk_comb} : {1'h0, p12_shifted_fraction};
  assign p13_rounded_fraction__1_comb = p13_do_round_up__6_comb ? {p13_add_8725_comb, p13_normal_chunk__1_comb} : {1'h0, p12_shifted_fraction__1};

  // Registers for pipe stage 13:
  reg [7:0] p13_greater_exp_bexp;
  reg [7:0] p13_greater_exp_bexp__1;
  reg [4:0] p13_encode_8552;
  reg [4:0] p13_encode_8553;
  reg [27:0] p13_rounded_fraction;
  reg [27:0] p13_rounded_fraction__1;
  reg p13_ne_8486;
  reg p13_ne_8487;
  reg p13_nor_8416;
  reg p13_nor_8418;
  reg p13_is_result_nan__5;
  reg p13_is_operand_inf;
  reg p13_is_result_nan__6;
  reg p13_is_operand_inf__1;
  reg [22:0] p13_in0_r_fraction__6;
  reg [7:0] p13_in0_r_bexp__6;
  reg [22:0] p13_in0_i_fraction__6;
  reg [7:0] p13_in0_i_bexp__6;
  reg p13_result_sign__13;
  reg p13_result_sign__14;
  reg p13_in0_r_sign__2;
  reg p13_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p13_greater_exp_bexp <= p12_greater_exp_bexp;
    p13_greater_exp_bexp__1 <= p12_greater_exp_bexp__1;
    p13_encode_8552 <= p12_encode_8552;
    p13_encode_8553 <= p12_encode_8553;
    p13_rounded_fraction <= p13_rounded_fraction_comb;
    p13_rounded_fraction__1 <= p13_rounded_fraction__1_comb;
    p13_ne_8486 <= p12_ne_8486;
    p13_ne_8487 <= p12_ne_8487;
    p13_nor_8416 <= p12_nor_8416;
    p13_nor_8418 <= p12_nor_8418;
    p13_is_result_nan__5 <= p12_is_result_nan__5;
    p13_is_operand_inf <= p12_is_operand_inf;
    p13_is_result_nan__6 <= p12_is_result_nan__6;
    p13_is_operand_inf__1 <= p12_is_operand_inf__1;
    p13_in0_r_fraction__6 <= p12_in0_r_fraction__6;
    p13_in0_r_bexp__6 <= p12_in0_r_bexp__6;
    p13_in0_i_fraction__6 <= p12_in0_i_fraction__6;
    p13_in0_i_bexp__6 <= p12_in0_i_bexp__6;
    p13_result_sign__13 <= p12_result_sign__13;
    p13_result_sign__14 <= p12_result_sign__14;
    p13_in0_r_sign__2 <= p12_in0_r_sign__2;
    p13_in0_i_sign__2 <= p12_in0_i_sign__2;
  end

  // ===== Pipe stage 14:
  wire p14_rounding_carry_comb;
  wire p14_rounding_carry__1_comb;
  wire [8:0] p14_add_8789_comb;
  wire [8:0] p14_add_8791_comb;
  wire [2:0] p14_add_8804_comb;
  wire [2:0] p14_add_8805_comb;
  wire [27:0] p14_shrl_8806_comb;
  wire [27:0] p14_shrl_8807_comb;
  wire [9:0] p14_add_8796_comb;
  wire [9:0] p14_add_8797_comb;
  wire [22:0] p14_result_fraction__13_comb;
  wire [22:0] p14_result_fraction__15_comb;
  assign p14_rounding_carry_comb = p13_rounded_fraction[27];
  assign p14_rounding_carry__1_comb = p13_rounded_fraction__1[27];
  assign p14_add_8789_comb = {1'h0, p13_greater_exp_bexp} + {8'h00, p14_rounding_carry_comb};
  assign p14_add_8791_comb = {1'h0, p13_greater_exp_bexp__1} + {8'h00, p14_rounding_carry__1_comb};
  assign p14_add_8804_comb = {2'h0, p14_rounding_carry_comb} + 3'h3;
  assign p14_add_8805_comb = {2'h0, p14_rounding_carry__1_comb} + 3'h3;
  assign p14_shrl_8806_comb = p13_rounded_fraction >> p14_add_8804_comb;
  assign p14_shrl_8807_comb = p13_rounded_fraction__1 >> p14_add_8805_comb;
  assign p14_add_8796_comb = {1'h0, p14_add_8789_comb} + 10'h001;
  assign p14_add_8797_comb = {1'h0, p14_add_8791_comb} + 10'h001;
  assign p14_result_fraction__13_comb = p14_shrl_8806_comb[22:0];
  assign p14_result_fraction__15_comb = p14_shrl_8807_comb[22:0];

  // Registers for pipe stage 14:
  reg [4:0] p14_encode_8552;
  reg [4:0] p14_encode_8553;
  reg [9:0] p14_add_8796;
  reg p14_ne_8486;
  reg [9:0] p14_add_8797;
  reg p14_ne_8487;
  reg p14_nor_8416;
  reg p14_nor_8418;
  reg [22:0] p14_result_fraction__13;
  reg p14_is_result_nan__5;
  reg p14_is_operand_inf;
  reg [22:0] p14_result_fraction__15;
  reg p14_is_result_nan__6;
  reg p14_is_operand_inf__1;
  reg [22:0] p14_in0_r_fraction__6;
  reg [7:0] p14_in0_r_bexp__6;
  reg [22:0] p14_in0_i_fraction__6;
  reg [7:0] p14_in0_i_bexp__6;
  reg p14_result_sign__13;
  reg p14_result_sign__14;
  reg p14_in0_r_sign__2;
  reg p14_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p14_encode_8552 <= p13_encode_8552;
    p14_encode_8553 <= p13_encode_8553;
    p14_add_8796 <= p14_add_8796_comb;
    p14_ne_8486 <= p13_ne_8486;
    p14_add_8797 <= p14_add_8797_comb;
    p14_ne_8487 <= p13_ne_8487;
    p14_nor_8416 <= p13_nor_8416;
    p14_nor_8418 <= p13_nor_8418;
    p14_result_fraction__13 <= p14_result_fraction__13_comb;
    p14_is_result_nan__5 <= p13_is_result_nan__5;
    p14_is_operand_inf <= p13_is_operand_inf;
    p14_result_fraction__15 <= p14_result_fraction__15_comb;
    p14_is_result_nan__6 <= p13_is_result_nan__6;
    p14_is_operand_inf__1 <= p13_is_operand_inf__1;
    p14_in0_r_fraction__6 <= p13_in0_r_fraction__6;
    p14_in0_r_bexp__6 <= p13_in0_r_bexp__6;
    p14_in0_i_fraction__6 <= p13_in0_i_fraction__6;
    p14_in0_i_bexp__6 <= p13_in0_i_bexp__6;
    p14_result_sign__13 <= p13_result_sign__13;
    p14_result_sign__14 <= p13_result_sign__14;
    p14_in0_r_sign__2 <= p13_in0_r_sign__2;
    p14_in0_i_sign__2 <= p13_in0_i_sign__2;
  end

  // ===== Pipe stage 15:
  wire [9:0] p15_wide_exponent_comb;
  wire [9:0] p15_wide_exponent__3_comb;
  wire [9:0] p15_wide_exponent__1_comb;
  wire [9:0] p15_wide_exponent__4_comb;
  wire p15_bit_slice_8864_comb;
  wire p15_bit_slice_8865_comb;
  wire [8:0] p15_bit_slice_8866_comb;
  wire [8:0] p15_bit_slice_8867_comb;
  assign p15_wide_exponent_comb = p14_add_8796 - {5'h00, p14_encode_8552};
  assign p15_wide_exponent__3_comb = p14_add_8797 - {5'h00, p14_encode_8553};
  assign p15_wide_exponent__1_comb = p15_wide_exponent_comb & {10{p14_ne_8486}};
  assign p15_wide_exponent__4_comb = p15_wide_exponent__3_comb & {10{p14_ne_8487}};
  assign p15_bit_slice_8864_comb = p15_wide_exponent__1_comb[9];
  assign p15_bit_slice_8865_comb = p15_wide_exponent__4_comb[9];
  assign p15_bit_slice_8866_comb = p15_wide_exponent__1_comb[8:0];
  assign p15_bit_slice_8867_comb = p15_wide_exponent__4_comb[8:0];

  // Registers for pipe stage 15:
  reg p15_bit_slice_8864;
  reg p15_bit_slice_8865;
  reg [8:0] p15_bit_slice_8866;
  reg [8:0] p15_bit_slice_8867;
  reg p15_nor_8416;
  reg p15_nor_8418;
  reg [22:0] p15_result_fraction__13;
  reg p15_is_result_nan__5;
  reg p15_is_operand_inf;
  reg [22:0] p15_result_fraction__15;
  reg p15_is_result_nan__6;
  reg p15_is_operand_inf__1;
  reg [22:0] p15_in0_r_fraction__6;
  reg [7:0] p15_in0_r_bexp__6;
  reg [22:0] p15_in0_i_fraction__6;
  reg [7:0] p15_in0_i_bexp__6;
  reg p15_result_sign__13;
  reg p15_result_sign__14;
  reg p15_in0_r_sign__2;
  reg p15_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p15_bit_slice_8864 <= p15_bit_slice_8864_comb;
    p15_bit_slice_8865 <= p15_bit_slice_8865_comb;
    p15_bit_slice_8866 <= p15_bit_slice_8866_comb;
    p15_bit_slice_8867 <= p15_bit_slice_8867_comb;
    p15_nor_8416 <= p14_nor_8416;
    p15_nor_8418 <= p14_nor_8418;
    p15_result_fraction__13 <= p14_result_fraction__13;
    p15_is_result_nan__5 <= p14_is_result_nan__5;
    p15_is_operand_inf <= p14_is_operand_inf;
    p15_result_fraction__15 <= p14_result_fraction__15;
    p15_is_result_nan__6 <= p14_is_result_nan__6;
    p15_is_operand_inf__1 <= p14_is_operand_inf__1;
    p15_in0_r_fraction__6 <= p14_in0_r_fraction__6;
    p15_in0_r_bexp__6 <= p14_in0_r_bexp__6;
    p15_in0_i_fraction__6 <= p14_in0_i_fraction__6;
    p15_in0_i_bexp__6 <= p14_in0_i_bexp__6;
    p15_result_sign__13 <= p14_result_sign__13;
    p15_result_sign__14 <= p14_result_sign__14;
    p15_in0_r_sign__2 <= p14_in0_r_sign__2;
    p15_in0_i_sign__2 <= p14_in0_i_sign__2;
  end

  // ===== Pipe stage 16:
  wire [8:0] p16_wide_exponent__2_comb;
  wire [8:0] p16_wide_exponent__5_comb;
  wire p16_bit_slice_8921_comb;
  wire p16_bit_slice_8929_comb;
  wire p16_bit_slice_8931_comb;
  wire p16_bit_slice_8933_comb;
  wire p16_or_8930_comb;
  wire p16_or_8932_comb;
  wire p16_and_8934_comb;
  wire p16_and_8935_comb;
  wire [7:0] p16_bit_slice_8936_comb;
  wire [7:0] p16_bit_slice_8937_comb;
  assign p16_wide_exponent__2_comb = p15_bit_slice_8866 & {9{~p15_bit_slice_8864}};
  assign p16_wide_exponent__5_comb = p15_bit_slice_8867 & {9{~p15_bit_slice_8865}};
  assign p16_bit_slice_8921_comb = p16_wide_exponent__2_comb[8];
  assign p16_bit_slice_8929_comb = p16_wide_exponent__5_comb[8];
  assign p16_bit_slice_8931_comb = p16_wide_exponent__2_comb[0];
  assign p16_bit_slice_8933_comb = p16_wide_exponent__5_comb[0];
  assign p16_or_8930_comb = p16_wide_exponent__2_comb[1] | p16_wide_exponent__2_comb[2] | p16_wide_exponent__2_comb[3] | p16_wide_exponent__2_comb[4] | p16_wide_exponent__2_comb[5] | p16_wide_exponent__2_comb[6] | p16_wide_exponent__2_comb[7] | p16_bit_slice_8921_comb;
  assign p16_or_8932_comb = p16_wide_exponent__5_comb[1] | p16_wide_exponent__5_comb[2] | p16_wide_exponent__5_comb[3] | p16_wide_exponent__5_comb[4] | p16_wide_exponent__5_comb[5] | p16_wide_exponent__5_comb[6] | p16_wide_exponent__5_comb[7] | p16_bit_slice_8929_comb;
  assign p16_and_8934_comb = p16_bit_slice_8931_comb & p16_wide_exponent__2_comb[1] & p16_wide_exponent__2_comb[2] & p16_wide_exponent__2_comb[3] & p16_wide_exponent__2_comb[4] & p16_wide_exponent__2_comb[5] & p16_wide_exponent__2_comb[6] & p16_wide_exponent__2_comb[7];
  assign p16_and_8935_comb = p16_bit_slice_8933_comb & p16_wide_exponent__5_comb[1] & p16_wide_exponent__5_comb[2] & p16_wide_exponent__5_comb[3] & p16_wide_exponent__5_comb[4] & p16_wide_exponent__5_comb[5] & p16_wide_exponent__5_comb[6] & p16_wide_exponent__5_comb[7];
  assign p16_bit_slice_8936_comb = p16_wide_exponent__2_comb[7:0];
  assign p16_bit_slice_8937_comb = p16_wide_exponent__5_comb[7:0];

  // Registers for pipe stage 16:
  reg p16_bit_slice_8921;
  reg p16_bit_slice_8929;
  reg p16_or_8930;
  reg p16_bit_slice_8931;
  reg p16_or_8932;
  reg p16_bit_slice_8933;
  reg p16_and_8934;
  reg p16_and_8935;
  reg p16_nor_8416;
  reg p16_nor_8418;
  reg [22:0] p16_result_fraction__13;
  reg p16_is_result_nan__5;
  reg p16_is_operand_inf;
  reg [22:0] p16_result_fraction__15;
  reg p16_is_result_nan__6;
  reg p16_is_operand_inf__1;
  reg [7:0] p16_bit_slice_8936;
  reg [7:0] p16_bit_slice_8937;
  reg [22:0] p16_in0_r_fraction__6;
  reg [7:0] p16_in0_r_bexp__6;
  reg [22:0] p16_in0_i_fraction__6;
  reg [7:0] p16_in0_i_bexp__6;
  reg p16_result_sign__13;
  reg p16_result_sign__14;
  reg p16_in0_r_sign__2;
  reg p16_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p16_bit_slice_8921 <= p16_bit_slice_8921_comb;
    p16_bit_slice_8929 <= p16_bit_slice_8929_comb;
    p16_or_8930 <= p16_or_8930_comb;
    p16_bit_slice_8931 <= p16_bit_slice_8931_comb;
    p16_or_8932 <= p16_or_8932_comb;
    p16_bit_slice_8933 <= p16_bit_slice_8933_comb;
    p16_and_8934 <= p16_and_8934_comb;
    p16_and_8935 <= p16_and_8935_comb;
    p16_nor_8416 <= p15_nor_8416;
    p16_nor_8418 <= p15_nor_8418;
    p16_result_fraction__13 <= p15_result_fraction__13;
    p16_is_result_nan__5 <= p15_is_result_nan__5;
    p16_is_operand_inf <= p15_is_operand_inf;
    p16_result_fraction__15 <= p15_result_fraction__15;
    p16_is_result_nan__6 <= p15_is_result_nan__6;
    p16_is_operand_inf__1 <= p15_is_operand_inf__1;
    p16_bit_slice_8936 <= p16_bit_slice_8936_comb;
    p16_bit_slice_8937 <= p16_bit_slice_8937_comb;
    p16_in0_r_fraction__6 <= p15_in0_r_fraction__6;
    p16_in0_r_bexp__6 <= p15_in0_r_bexp__6;
    p16_in0_i_fraction__6 <= p15_in0_i_fraction__6;
    p16_in0_i_bexp__6 <= p15_in0_i_bexp__6;
    p16_result_sign__13 <= p15_result_sign__13;
    p16_result_sign__14 <= p15_result_sign__14;
    p16_in0_r_sign__2 <= p15_in0_r_sign__2;
    p16_in0_i_sign__2 <= p15_in0_i_sign__2;
  end

  // ===== Pipe stage 17:
  wire p17_nor_8993_comb;
  wire p17_nor_8995_comb;
  wire [22:0] p17_result_fraction__14_comb;
  wire [22:0] p17_nan_fraction__14_comb;
  wire [7:0] p17_high_exp__36_comb;
  wire [22:0] p17_result_fraction__16_comb;
  wire [22:0] p17_nan_fraction__15_comb;
  wire [7:0] p17_high_exp__37_comb;
  wire [22:0] p17_result_fraction__17_comb;
  wire [7:0] p17_result_exponent__2_comb;
  wire [22:0] p17_result_fraction__18_comb;
  wire [7:0] p17_result_exponent__1_comb;
  assign p17_nor_8993_comb = ~(p16_bit_slice_8921 | p16_and_8934);
  assign p17_nor_8995_comb = ~(p16_bit_slice_8929 | p16_and_8935);
  assign p17_result_fraction__14_comb = p16_result_fraction__13 & {23{~(~(p16_or_8930 | p16_bit_slice_8931))}} & {23{p17_nor_8993_comb}} & {23{p16_nor_8416}};
  assign p17_nan_fraction__14_comb = 23'h40_0000;
  assign p17_high_exp__36_comb = 8'hff;
  assign p17_result_fraction__16_comb = p16_result_fraction__15 & {23{~(~(p16_or_8932 | p16_bit_slice_8933))}} & {23{p17_nor_8995_comb}} & {23{p16_nor_8418}};
  assign p17_nan_fraction__15_comb = 23'h40_0000;
  assign p17_high_exp__37_comb = 8'hff;
  assign p17_result_fraction__17_comb = p16_is_result_nan__5 ? p17_nan_fraction__14_comb : p17_result_fraction__14_comb;
  assign p17_result_exponent__2_comb = p16_is_result_nan__5 | p16_is_operand_inf | ~p17_nor_8993_comb ? p17_high_exp__36_comb : p16_bit_slice_8936;
  assign p17_result_fraction__18_comb = p16_is_result_nan__6 ? p17_nan_fraction__15_comb : p17_result_fraction__16_comb;
  assign p17_result_exponent__1_comb = p16_is_result_nan__6 | p16_is_operand_inf__1 | ~p17_nor_8995_comb ? p17_high_exp__37_comb : p16_bit_slice_8937;

  // Registers for pipe stage 17:
  reg [22:0] p17_in0_r_fraction__6;
  reg [7:0] p17_in0_r_bexp__6;
  reg [22:0] p17_result_fraction__17;
  reg [7:0] p17_result_exponent__2;
  reg [22:0] p17_in0_i_fraction__6;
  reg [7:0] p17_in0_i_bexp__6;
  reg [22:0] p17_result_fraction__18;
  reg [7:0] p17_result_exponent__1;
  reg p17_result_sign__13;
  reg p17_result_sign__14;
  reg p17_in0_r_sign__2;
  reg p17_in0_i_sign__2;
  always_ff @ (posedge clk) begin
    p17_in0_r_fraction__6 <= p16_in0_r_fraction__6;
    p17_in0_r_bexp__6 <= p16_in0_r_bexp__6;
    p17_result_fraction__17 <= p17_result_fraction__17_comb;
    p17_result_exponent__2 <= p17_result_exponent__2_comb;
    p17_in0_i_fraction__6 <= p16_in0_i_fraction__6;
    p17_in0_i_bexp__6 <= p16_in0_i_bexp__6;
    p17_result_fraction__18 <= p17_result_fraction__18_comb;
    p17_result_exponent__1 <= p17_result_exponent__1_comb;
    p17_result_sign__13 <= p16_result_sign__13;
    p17_result_sign__14 <= p16_result_sign__14;
    p17_in0_r_sign__2 <= p16_in0_r_sign__2;
    p17_in0_i_sign__2 <= p16_in0_i_sign__2;
  end

  // ===== Pipe stage 18:
  wire [5:0] p18_add_9067_comb;
  wire p18_ugt_9069_comb;
  wire [5:0] p18_add_9073_comb;
  wire [5:0] p18_add_9078_comb;
  wire p18_ugt_9080_comb;
  wire [5:0] p18_add_9084_comb;
  wire [27:0] p18_wide_x__4_comb;
  wire [7:0] p18_greater_exp_bexp__2_comb;
  wire [27:0] p18_wide_y__4_comb;
  wire [27:0] p18_wide_x__6_comb;
  wire [7:0] p18_greater_exp_bexp__3_comb;
  wire [27:0] p18_wide_y__6_comb;
  wire [27:0] p18_wide_x__5_comb;
  wire [7:0] p18_sub_9101_comb;
  wire [27:0] p18_wide_y__5_comb;
  wire [7:0] p18_sub_9103_comb;
  wire [27:0] p18_wide_x__7_comb;
  wire [7:0] p18_sub_9105_comb;
  wire [27:0] p18_wide_y__7_comb;
  wire [7:0] p18_sub_9107_comb;
  wire p18_eq_9111_comb;
  wire p18_eq_9114_comb;
  wire p18_ne_9116_comb;
  wire p18_eq_9117_comb;
  wire p18_ne_9118_comb;
  wire p18_eq_9119_comb;
  wire p18_ne_9122_comb;
  wire p18_ne_9123_comb;
  assign p18_add_9067_comb = p17_in0_r_bexp__6[7:2] + 6'h07;
  assign p18_ugt_9069_comb = p17_in0_r_bexp__6 > p17_result_exponent__2;
  assign p18_add_9073_comb = p17_result_exponent__2[7:2] + 6'h07;
  assign p18_add_9078_comb = p17_in0_i_bexp__6[7:2] + 6'h07;
  assign p18_ugt_9080_comb = p17_in0_i_bexp__6 > p17_result_exponent__1;
  assign p18_add_9084_comb = p17_result_exponent__1[7:2] + 6'h07;
  assign p18_wide_x__4_comb = {{2'h0, p17_in0_r_fraction__6} | 25'h080_0000, 3'h0};
  assign p18_greater_exp_bexp__2_comb = p18_ugt_9069_comb ? p17_in0_r_bexp__6 : p17_result_exponent__2;
  assign p18_wide_y__4_comb = {{2'h0, p17_result_fraction__17} | 25'h080_0000, 3'h0};
  assign p18_wide_x__6_comb = {{2'h0, p17_in0_i_fraction__6} | 25'h080_0000, 3'h0};
  assign p18_greater_exp_bexp__3_comb = p18_ugt_9080_comb ? p17_in0_i_bexp__6 : p17_result_exponent__1;
  assign p18_wide_y__6_comb = {{2'h0, p17_result_fraction__18} | 25'h080_0000, 3'h0};
  assign p18_wide_x__5_comb = p18_wide_x__4_comb & {28{p17_in0_r_bexp__6 != 8'h00}};
  assign p18_sub_9101_comb = {p18_add_9067_comb, p17_in0_r_bexp__6[1:0]} - p18_greater_exp_bexp__2_comb;
  assign p18_wide_y__5_comb = p18_wide_y__4_comb & {28{p17_result_exponent__2 != 8'h00}};
  assign p18_sub_9103_comb = {p18_add_9073_comb, p17_result_exponent__2[1:0]} - p18_greater_exp_bexp__2_comb;
  assign p18_wide_x__7_comb = p18_wide_x__6_comb & {28{p17_in0_i_bexp__6 != 8'h00}};
  assign p18_sub_9105_comb = {p18_add_9078_comb, p17_in0_i_bexp__6[1:0]} - p18_greater_exp_bexp__3_comb;
  assign p18_wide_y__7_comb = p18_wide_y__6_comb & {28{p17_result_exponent__1 != 8'h00}};
  assign p18_sub_9107_comb = {p18_add_9084_comb, p17_result_exponent__1[1:0]} - p18_greater_exp_bexp__3_comb;
  assign p18_eq_9111_comb = p17_result_fraction__17 == 23'h00_0000;
  assign p18_eq_9114_comb = p17_result_fraction__18 == 23'h00_0000;
  assign p18_ne_9116_comb = p17_in0_r_fraction__6 != 23'h00_0000;
  assign p18_eq_9117_comb = p17_in0_r_fraction__6 == 23'h00_0000;
  assign p18_ne_9118_comb = p17_in0_i_fraction__6 != 23'h00_0000;
  assign p18_eq_9119_comb = p17_in0_i_fraction__6 == 23'h00_0000;
  assign p18_ne_9122_comb = p17_result_fraction__17 != 23'h00_0000;
  assign p18_ne_9123_comb = p17_result_fraction__18 != 23'h00_0000;

  // Registers for pipe stage 18:
  reg [7:0] p18_in0_r_bexp__6;
  reg [7:0] p18_result_exponent__2;
  reg [7:0] p18_in0_i_bexp__6;
  reg [7:0] p18_result_exponent__1;
  reg p18_ugt_9069;
  reg p18_ugt_9080;
  reg [7:0] p18_greater_exp_bexp__2;
  reg [7:0] p18_greater_exp_bexp__3;
  reg [27:0] p18_wide_x__5;
  reg [7:0] p18_sub_9101;
  reg [27:0] p18_wide_y__5;
  reg [7:0] p18_sub_9103;
  reg [27:0] p18_wide_x__7;
  reg [7:0] p18_sub_9105;
  reg [27:0] p18_wide_y__7;
  reg [7:0] p18_sub_9107;
  reg p18_result_sign__13;
  reg p18_result_sign__14;
  reg p18_in0_r_sign__2;
  reg p18_in0_i_sign__2;
  reg p18_eq_9111;
  reg p18_eq_9114;
  reg p18_ne_9116;
  reg p18_eq_9117;
  reg p18_ne_9118;
  reg p18_eq_9119;
  reg p18_ne_9122;
  reg p18_ne_9123;
  always_ff @ (posedge clk) begin
    p18_in0_r_bexp__6 <= p17_in0_r_bexp__6;
    p18_result_exponent__2 <= p17_result_exponent__2;
    p18_in0_i_bexp__6 <= p17_in0_i_bexp__6;
    p18_result_exponent__1 <= p17_result_exponent__1;
    p18_ugt_9069 <= p18_ugt_9069_comb;
    p18_ugt_9080 <= p18_ugt_9080_comb;
    p18_greater_exp_bexp__2 <= p18_greater_exp_bexp__2_comb;
    p18_greater_exp_bexp__3 <= p18_greater_exp_bexp__3_comb;
    p18_wide_x__5 <= p18_wide_x__5_comb;
    p18_sub_9101 <= p18_sub_9101_comb;
    p18_wide_y__5 <= p18_wide_y__5_comb;
    p18_sub_9103 <= p18_sub_9103_comb;
    p18_wide_x__7 <= p18_wide_x__7_comb;
    p18_sub_9105 <= p18_sub_9105_comb;
    p18_wide_y__7 <= p18_wide_y__7_comb;
    p18_sub_9107 <= p18_sub_9107_comb;
    p18_result_sign__13 <= p17_result_sign__13;
    p18_result_sign__14 <= p17_result_sign__14;
    p18_in0_r_sign__2 <= p17_in0_r_sign__2;
    p18_in0_i_sign__2 <= p17_in0_i_sign__2;
    p18_eq_9111 <= p18_eq_9111_comb;
    p18_eq_9114 <= p18_eq_9114_comb;
    p18_ne_9116 <= p18_ne_9116_comb;
    p18_eq_9117 <= p18_eq_9117_comb;
    p18_ne_9118 <= p18_ne_9118_comb;
    p18_eq_9119 <= p18_eq_9119_comb;
    p18_ne_9122 <= p18_ne_9122_comb;
    p18_ne_9123 <= p18_ne_9123_comb;
  end

  // ===== Pipe stage 19:
  wire [27:0] p19_dropped_x__2_comb;
  wire [27:0] p19_dropped_y__2_comb;
  wire [27:0] p19_dropped_x__3_comb;
  wire [27:0] p19_dropped_y__3_comb;
  wire [7:0] p19_high_exp__38_comb;
  wire [7:0] p19_high_exp__39_comb;
  wire [7:0] p19_high_exp__40_comb;
  wire [7:0] p19_high_exp__41_comb;
  wire [7:0] p19_shift_x__2_comb;
  wire p19_sticky_x__2_comb;
  wire [7:0] p19_shift_y__2_comb;
  wire p19_sticky_y__2_comb;
  wire [7:0] p19_shift_x__3_comb;
  wire p19_sticky_x__3_comb;
  wire [7:0] p19_shift_y__3_comb;
  wire p19_sticky_y__3_comb;
  wire [7:0] p19_high_exp__46_comb;
  wire [7:0] p19_high_exp__47_comb;
  wire p19_eq_9228_comb;
  wire p19_eq_9221_comb;
  wire p19_eq_9231_comb;
  wire p19_eq_9224_comb;
  wire [27:0] p19_shifted_x__2_comb;
  wire [27:0] p19_shifted_y__2_comb;
  wire [27:0] p19_shifted_x__3_comb;
  wire [27:0] p19_shifted_y__3_comb;
  wire p19_and_9236_comb;
  wire p19_and_9237_comb;
  wire p19_and_9238_comb;
  wire p19_and_9239_comb;
  wire p19_re__1_sign_comb;
  wire p19_im__1_sign_comb;
  wire [27:0] p19_addend_x__4_comb;
  wire [27:0] p19_addend_y__4_comb;
  wire [27:0] p19_addend_x__6_comb;
  wire [27:0] p19_addend_y__6_comb;
  wire p19_nand_9227_comb;
  wire p19_nand_9230_comb;
  wire p19_nor_9232_comb;
  wire p19_and_9233_comb;
  wire p19_nor_9234_comb;
  wire p19_and_9235_comb;
  wire p19_and_9240_comb;
  wire p19_and_9241_comb;
  wire p19_nor_9242_comb;
  wire p19_and_9243_comb;
  wire p19_and_9244_comb;
  wire p19_nor_9245_comb;
  wire p19_is_operand_inf__2_comb;
  wire p19_is_operand_inf__3_comb;
  assign p19_dropped_x__2_comb = p18_sub_9101 >= 8'h1c ? 28'h000_0000 : p18_wide_x__5 << p18_sub_9101;
  assign p19_dropped_y__2_comb = p18_sub_9103 >= 8'h1c ? 28'h000_0000 : p18_wide_y__5 << p18_sub_9103;
  assign p19_dropped_x__3_comb = p18_sub_9105 >= 8'h1c ? 28'h000_0000 : p18_wide_x__7 << p18_sub_9105;
  assign p19_dropped_y__3_comb = p18_sub_9107 >= 8'h1c ? 28'h000_0000 : p18_wide_y__7 << p18_sub_9107;
  assign p19_high_exp__38_comb = 8'hff;
  assign p19_high_exp__39_comb = 8'hff;
  assign p19_high_exp__40_comb = 8'hff;
  assign p19_high_exp__41_comb = 8'hff;
  assign p19_shift_x__2_comb = p18_greater_exp_bexp__2 - p18_in0_r_bexp__6;
  assign p19_sticky_x__2_comb = p19_dropped_x__2_comb[27:3] != 25'h000_0000;
  assign p19_shift_y__2_comb = p18_greater_exp_bexp__2 - p18_result_exponent__2;
  assign p19_sticky_y__2_comb = p19_dropped_y__2_comb[27:3] != 25'h000_0000;
  assign p19_shift_x__3_comb = p18_greater_exp_bexp__3 - p18_in0_i_bexp__6;
  assign p19_sticky_x__3_comb = p19_dropped_x__3_comb[27:3] != 25'h000_0000;
  assign p19_shift_y__3_comb = p18_greater_exp_bexp__3 - p18_result_exponent__1;
  assign p19_sticky_y__3_comb = p19_dropped_y__3_comb[27:3] != 25'h000_0000;
  assign p19_high_exp__46_comb = 8'hff;
  assign p19_high_exp__47_comb = 8'hff;
  assign p19_eq_9228_comb = p18_in0_r_bexp__6 == p19_high_exp__38_comb;
  assign p19_eq_9221_comb = p18_result_exponent__2 == p19_high_exp__39_comb;
  assign p19_eq_9231_comb = p18_in0_i_bexp__6 == p19_high_exp__40_comb;
  assign p19_eq_9224_comb = p18_result_exponent__1 == p19_high_exp__41_comb;
  assign p19_shifted_x__2_comb = p19_shift_x__2_comb >= 8'h1c ? 28'h000_0000 : p18_wide_x__5 >> p19_shift_x__2_comb;
  assign p19_shifted_y__2_comb = p19_shift_y__2_comb >= 8'h1c ? 28'h000_0000 : p18_wide_y__5 >> p19_shift_y__2_comb;
  assign p19_shifted_x__3_comb = p19_shift_x__3_comb >= 8'h1c ? 28'h000_0000 : p18_wide_x__7 >> p19_shift_x__3_comb;
  assign p19_shifted_y__3_comb = p19_shift_y__3_comb >= 8'h1c ? 28'h000_0000 : p18_wide_y__7 >> p19_shift_y__3_comb;
  assign p19_and_9236_comb = p19_eq_9228_comb & p18_eq_9117;
  assign p19_and_9237_comb = p19_eq_9221_comb & p18_eq_9111;
  assign p19_and_9238_comb = p19_eq_9231_comb & p18_eq_9119;
  assign p19_and_9239_comb = p19_eq_9224_comb & p18_eq_9114;
  assign p19_re__1_sign_comb = ~p18_result_sign__13;
  assign p19_im__1_sign_comb = ~p18_result_sign__14;
  assign p19_addend_x__4_comb = p19_shifted_x__2_comb | {27'h000_0000, p19_sticky_x__2_comb};
  assign p19_addend_y__4_comb = p19_shifted_y__2_comb | {27'h000_0000, p19_sticky_y__2_comb};
  assign p19_addend_x__6_comb = p19_shifted_x__3_comb | {27'h000_0000, p19_sticky_x__3_comb};
  assign p19_addend_y__6_comb = p19_shifted_y__3_comb | {27'h000_0000, p19_sticky_y__3_comb};
  assign p19_nand_9227_comb = ~(p19_eq_9221_comb & p18_eq_9111);
  assign p19_nand_9230_comb = ~(p19_eq_9224_comb & p18_eq_9114);
  assign p19_nor_9232_comb = ~(p18_in0_r_bexp__6 != p19_high_exp__46_comb | p18_ne_9116 | p18_in0_r_sign__2);
  assign p19_and_9233_comb = p19_eq_9228_comb & p18_eq_9117 & p18_in0_r_sign__2;
  assign p19_nor_9234_comb = ~(p18_in0_i_bexp__6 != p19_high_exp__47_comb | p18_ne_9118 | p18_in0_i_sign__2);
  assign p19_and_9235_comb = p19_eq_9231_comb & p18_eq_9119 & p18_in0_i_sign__2;
  assign p19_and_9240_comb = p19_eq_9228_comb & p18_ne_9116;
  assign p19_and_9241_comb = p19_eq_9221_comb & p18_ne_9122;
  assign p19_nor_9242_comb = ~(p19_and_9236_comb | p19_and_9237_comb);
  assign p19_and_9243_comb = p19_eq_9231_comb & p18_ne_9118;
  assign p19_and_9244_comb = p19_eq_9224_comb & p18_ne_9123;
  assign p19_nor_9245_comb = ~(p19_and_9238_comb | p19_and_9239_comb);
  assign p19_is_operand_inf__2_comb = p19_and_9236_comb | p19_and_9237_comb;
  assign p19_is_operand_inf__3_comb = p19_and_9238_comb | p19_and_9239_comb;

  // Registers for pipe stage 19:
  reg p19_ugt_9069;
  reg p19_ugt_9080;
  reg [7:0] p19_greater_exp_bexp__2;
  reg [7:0] p19_greater_exp_bexp__3;
  reg p19_result_sign__13;
  reg p19_result_sign__14;
  reg p19_in0_r_sign__2;
  reg p19_in0_i_sign__2;
  reg p19_re__1_sign;
  reg p19_im__1_sign;
  reg [27:0] p19_addend_x__4;
  reg [27:0] p19_addend_y__4;
  reg [27:0] p19_addend_x__6;
  reg [27:0] p19_addend_y__6;
  reg p19_nand_9227;
  reg p19_nand_9230;
  reg p19_nor_9232;
  reg p19_and_9233;
  reg p19_nor_9234;
  reg p19_and_9235;
  reg p19_and_9240;
  reg p19_and_9241;
  reg p19_nor_9242;
  reg p19_and_9243;
  reg p19_and_9244;
  reg p19_nor_9245;
  reg p19_is_operand_inf__2;
  reg p19_is_operand_inf__3;
  always_ff @ (posedge clk) begin
    p19_ugt_9069 <= p18_ugt_9069;
    p19_ugt_9080 <= p18_ugt_9080;
    p19_greater_exp_bexp__2 <= p18_greater_exp_bexp__2;
    p19_greater_exp_bexp__3 <= p18_greater_exp_bexp__3;
    p19_result_sign__13 <= p18_result_sign__13;
    p19_result_sign__14 <= p18_result_sign__14;
    p19_in0_r_sign__2 <= p18_in0_r_sign__2;
    p19_in0_i_sign__2 <= p18_in0_i_sign__2;
    p19_re__1_sign <= p19_re__1_sign_comb;
    p19_im__1_sign <= p19_im__1_sign_comb;
    p19_addend_x__4 <= p19_addend_x__4_comb;
    p19_addend_y__4 <= p19_addend_y__4_comb;
    p19_addend_x__6 <= p19_addend_x__6_comb;
    p19_addend_y__6 <= p19_addend_y__6_comb;
    p19_nand_9227 <= p19_nand_9227_comb;
    p19_nand_9230 <= p19_nand_9230_comb;
    p19_nor_9232 <= p19_nor_9232_comb;
    p19_and_9233 <= p19_and_9233_comb;
    p19_nor_9234 <= p19_nor_9234_comb;
    p19_and_9235 <= p19_and_9235_comb;
    p19_and_9240 <= p19_and_9240_comb;
    p19_and_9241 <= p19_and_9241_comb;
    p19_nor_9242 <= p19_nor_9242_comb;
    p19_and_9243 <= p19_and_9243_comb;
    p19_and_9244 <= p19_and_9244_comb;
    p19_nor_9245 <= p19_nor_9245_comb;
    p19_is_operand_inf__2 <= p19_is_operand_inf__2_comb;
    p19_is_operand_inf__3 <= p19_is_operand_inf__3_comb;
  end

  // ===== Pipe stage 20:
  wire p20_greater_exp_sign__2_comb;
  wire p20_greater_exp_sign__3_comb;
  wire p20_greater_exp_sign__4_comb;
  wire p20_greater_exp_sign__5_comb;
  wire p20_nor_9340_comb;
  wire p20_nor_9341_comb;
  wire p20_nor_9342_comb;
  wire p20_nor_9343_comb;
  wire [27:0] p20_addend_x__5_comb;
  wire [27:0] p20_addend_y__5_comb;
  wire [27:0] p20_addend_x__7_comb;
  wire [27:0] p20_addend_y__7_comb;
  wire [27:0] p20_addend_x__9_comb;
  wire [27:0] p20_addend_y__9_comb;
  wire [27:0] p20_addend_x__11_comb;
  wire [27:0] p20_addend_y__11_comb;
  wire p20_has_pos_inf__2_comb;
  wire p20_has_neg_inf__2_comb;
  wire p20_has_pos_inf__3_comb;
  wire p20_has_neg_inf__3_comb;
  wire p20_has_pos_inf__4_comb;
  wire p20_has_neg_inf__4_comb;
  wire p20_has_pos_inf__5_comb;
  wire p20_has_neg_inf__5_comb;
  wire [28:0] p20_fraction__35_comb;
  wire [28:0] p20_fraction__36_comb;
  wire [28:0] p20_fraction__37_comb;
  wire [28:0] p20_fraction__38_comb;
  wire p20_is_result_nan__7_comb;
  wire p20_not_9357_comb;
  wire p20_is_result_nan__8_comb;
  wire p20_not_9359_comb;
  wire p20_is_result_nan__9_comb;
  wire p20_not_9361_comb;
  wire p20_is_result_nan__10_comb;
  wire p20_not_9363_comb;
  assign p20_greater_exp_sign__2_comb = p19_ugt_9069 ? p19_in0_r_sign__2 : p19_result_sign__13;
  assign p20_greater_exp_sign__3_comb = p19_ugt_9080 ? p19_in0_i_sign__2 : p19_result_sign__14;
  assign p20_greater_exp_sign__4_comb = p19_ugt_9069 ? p19_in0_r_sign__2 : p19_re__1_sign;
  assign p20_greater_exp_sign__5_comb = p19_ugt_9080 ? p19_in0_i_sign__2 : p19_im__1_sign;
  assign p20_nor_9340_comb = ~(p19_nand_9227 | p19_result_sign__13);
  assign p20_nor_9341_comb = ~(p19_nand_9227 | p19_re__1_sign);
  assign p20_nor_9342_comb = ~(p19_nand_9230 | p19_result_sign__14);
  assign p20_nor_9343_comb = ~(p19_nand_9230 | p19_im__1_sign);
  assign p20_addend_x__5_comb = p19_in0_r_sign__2 ^ p20_greater_exp_sign__2_comb ? -p19_addend_x__4 : p19_addend_x__4;
  assign p20_addend_y__5_comb = p19_result_sign__13 ^ p20_greater_exp_sign__2_comb ? -p19_addend_y__4 : p19_addend_y__4;
  assign p20_addend_x__7_comb = p19_in0_i_sign__2 ^ p20_greater_exp_sign__3_comb ? -p19_addend_x__6 : p19_addend_x__6;
  assign p20_addend_y__7_comb = p19_result_sign__14 ^ p20_greater_exp_sign__3_comb ? -p19_addend_y__6 : p19_addend_y__6;
  assign p20_addend_x__9_comb = p19_in0_r_sign__2 ^ p20_greater_exp_sign__4_comb ? -p19_addend_x__4 : p19_addend_x__4;
  assign p20_addend_y__9_comb = p19_re__1_sign ^ p20_greater_exp_sign__4_comb ? -p19_addend_y__4 : p19_addend_y__4;
  assign p20_addend_x__11_comb = p19_in0_i_sign__2 ^ p20_greater_exp_sign__5_comb ? -p19_addend_x__6 : p19_addend_x__6;
  assign p20_addend_y__11_comb = p19_im__1_sign ^ p20_greater_exp_sign__5_comb ? -p19_addend_y__6 : p19_addend_y__6;
  assign p20_has_pos_inf__2_comb = p19_nor_9232 | p20_nor_9340_comb;
  assign p20_has_neg_inf__2_comb = p19_and_9233 | p20_nor_9341_comb;
  assign p20_has_pos_inf__3_comb = p19_nor_9234 | p20_nor_9342_comb;
  assign p20_has_neg_inf__3_comb = p19_and_9235 | p20_nor_9343_comb;
  assign p20_has_pos_inf__4_comb = p19_nor_9232 | p20_nor_9341_comb;
  assign p20_has_neg_inf__4_comb = p19_and_9233 | p20_nor_9340_comb;
  assign p20_has_pos_inf__5_comb = p19_nor_9234 | p20_nor_9343_comb;
  assign p20_has_neg_inf__5_comb = p19_and_9235 | p20_nor_9342_comb;
  assign p20_fraction__35_comb = {{1{p20_addend_x__5_comb[27]}}, p20_addend_x__5_comb} + {{1{p20_addend_y__5_comb[27]}}, p20_addend_y__5_comb};
  assign p20_fraction__36_comb = {{1{p20_addend_x__7_comb[27]}}, p20_addend_x__7_comb} + {{1{p20_addend_y__7_comb[27]}}, p20_addend_y__7_comb};
  assign p20_fraction__37_comb = {{1{p20_addend_x__9_comb[27]}}, p20_addend_x__9_comb} + {{1{p20_addend_y__9_comb[27]}}, p20_addend_y__9_comb};
  assign p20_fraction__38_comb = {{1{p20_addend_x__11_comb[27]}}, p20_addend_x__11_comb} + {{1{p20_addend_y__11_comb[27]}}, p20_addend_y__11_comb};
  assign p20_is_result_nan__7_comb = p19_and_9240 | p19_and_9241 | p20_has_pos_inf__2_comb & p20_has_neg_inf__2_comb;
  assign p20_not_9357_comb = ~p20_has_pos_inf__2_comb;
  assign p20_is_result_nan__8_comb = p19_and_9243 | p19_and_9244 | p20_has_pos_inf__3_comb & p20_has_neg_inf__3_comb;
  assign p20_not_9359_comb = ~p20_has_pos_inf__3_comb;
  assign p20_is_result_nan__9_comb = p19_and_9240 | p19_and_9241 | p20_has_pos_inf__4_comb & p20_has_neg_inf__4_comb;
  assign p20_not_9361_comb = ~p20_has_pos_inf__4_comb;
  assign p20_is_result_nan__10_comb = p19_and_9243 | p19_and_9244 | p20_has_pos_inf__5_comb & p20_has_neg_inf__5_comb;
  assign p20_not_9363_comb = ~p20_has_pos_inf__5_comb;

  // Registers for pipe stage 20:
  reg [7:0] p20_greater_exp_bexp__2;
  reg [7:0] p20_greater_exp_bexp__3;
  reg p20_greater_exp_sign__2;
  reg p20_greater_exp_sign__3;
  reg p20_greater_exp_sign__4;
  reg p20_greater_exp_sign__5;
  reg [28:0] p20_fraction__35;
  reg [28:0] p20_fraction__36;
  reg [28:0] p20_fraction__37;
  reg [28:0] p20_fraction__38;
  reg p20_nor_9242;
  reg p20_nor_9245;
  reg p20_is_result_nan__7;
  reg p20_is_operand_inf__2;
  reg p20_not_9357;
  reg p20_is_result_nan__8;
  reg p20_is_operand_inf__3;
  reg p20_not_9359;
  reg p20_is_result_nan__9;
  reg p20_not_9361;
  reg p20_is_result_nan__10;
  reg p20_not_9363;
  always_ff @ (posedge clk) begin
    p20_greater_exp_bexp__2 <= p19_greater_exp_bexp__2;
    p20_greater_exp_bexp__3 <= p19_greater_exp_bexp__3;
    p20_greater_exp_sign__2 <= p20_greater_exp_sign__2_comb;
    p20_greater_exp_sign__3 <= p20_greater_exp_sign__3_comb;
    p20_greater_exp_sign__4 <= p20_greater_exp_sign__4_comb;
    p20_greater_exp_sign__5 <= p20_greater_exp_sign__5_comb;
    p20_fraction__35 <= p20_fraction__35_comb;
    p20_fraction__36 <= p20_fraction__36_comb;
    p20_fraction__37 <= p20_fraction__37_comb;
    p20_fraction__38 <= p20_fraction__38_comb;
    p20_nor_9242 <= p19_nor_9242;
    p20_nor_9245 <= p19_nor_9245;
    p20_is_result_nan__7 <= p20_is_result_nan__7_comb;
    p20_is_operand_inf__2 <= p19_is_operand_inf__2;
    p20_not_9357 <= p20_not_9357_comb;
    p20_is_result_nan__8 <= p20_is_result_nan__8_comb;
    p20_is_operand_inf__3 <= p19_is_operand_inf__3;
    p20_not_9359 <= p20_not_9359_comb;
    p20_is_result_nan__9 <= p20_is_result_nan__9_comb;
    p20_not_9361 <= p20_not_9361_comb;
    p20_is_result_nan__10 <= p20_is_result_nan__10_comb;
    p20_not_9363 <= p20_not_9363_comb;
  end

  // ===== Pipe stage 21:
  wire p21_fraction_is_zero__2_comb;
  wire p21_fraction_is_zero__3_comb;
  wire p21_fraction_is_zero__4_comb;
  wire p21_fraction_is_zero__5_comb;
  wire p21_result_sign__15_comb;
  wire p21_result_sign__17_comb;
  wire p21_result_sign__20_comb;
  wire p21_result_sign__23_comb;
  wire [27:0] p21_abs_fraction__2_comb;
  wire [27:0] p21_abs_fraction__3_comb;
  wire [27:0] p21_abs_fraction__4_comb;
  wire [27:0] p21_abs_fraction__5_comb;
  wire p21_ne_9428_comb;
  wire p21_ne_9429_comb;
  wire p21_ne_9430_comb;
  wire p21_ne_9431_comb;
  wire p21_result_sign__16_comb;
  wire p21_result_sign__18_comb;
  wire p21_result_sign__21_comb;
  wire p21_result_sign__24_comb;
  assign p21_fraction_is_zero__2_comb = p20_fraction__35 == 29'h0000_0000;
  assign p21_fraction_is_zero__3_comb = p20_fraction__36 == 29'h0000_0000;
  assign p21_fraction_is_zero__4_comb = p20_fraction__37 == 29'h0000_0000;
  assign p21_fraction_is_zero__5_comb = p20_fraction__38 == 29'h0000_0000;
  assign p21_result_sign__15_comb = ~(~p20_fraction__35[28] | p20_greater_exp_sign__2) | ~(p20_fraction__35[28] | p21_fraction_is_zero__2_comb | ~p20_greater_exp_sign__2);
  assign p21_result_sign__17_comb = ~(~p20_fraction__36[28] | p20_greater_exp_sign__3) | ~(p20_fraction__36[28] | p21_fraction_is_zero__3_comb | ~p20_greater_exp_sign__3);
  assign p21_result_sign__20_comb = ~(~p20_fraction__37[28] | p20_greater_exp_sign__4) | ~(p20_fraction__37[28] | p21_fraction_is_zero__4_comb | ~p20_greater_exp_sign__4);
  assign p21_result_sign__23_comb = ~(~p20_fraction__38[28] | p20_greater_exp_sign__5) | ~(p20_fraction__38[28] | p21_fraction_is_zero__5_comb | ~p20_greater_exp_sign__5);
  assign p21_abs_fraction__2_comb = p20_fraction__35[28] ? -p20_fraction__35[27:0] : p20_fraction__35[27:0];
  assign p21_abs_fraction__3_comb = p20_fraction__36[28] ? -p20_fraction__36[27:0] : p20_fraction__36[27:0];
  assign p21_abs_fraction__4_comb = p20_fraction__37[28] ? -p20_fraction__37[27:0] : p20_fraction__37[27:0];
  assign p21_abs_fraction__5_comb = p20_fraction__38[28] ? -p20_fraction__38[27:0] : p20_fraction__38[27:0];
  assign p21_ne_9428_comb = p20_fraction__35 != 29'h0000_0000;
  assign p21_ne_9429_comb = p20_fraction__36 != 29'h0000_0000;
  assign p21_ne_9430_comb = p20_fraction__37 != 29'h0000_0000;
  assign p21_ne_9431_comb = p20_fraction__38 != 29'h0000_0000;
  assign p21_result_sign__16_comb = p20_is_operand_inf__2 ? p20_not_9357 : p21_result_sign__15_comb;
  assign p21_result_sign__18_comb = p20_is_operand_inf__3 ? p20_not_9359 : p21_result_sign__17_comb;
  assign p21_result_sign__21_comb = p20_is_operand_inf__2 ? p20_not_9361 : p21_result_sign__20_comb;
  assign p21_result_sign__24_comb = p20_is_operand_inf__3 ? p20_not_9363 : p21_result_sign__23_comb;

  // Registers for pipe stage 21:
  reg [7:0] p21_greater_exp_bexp__2;
  reg [7:0] p21_greater_exp_bexp__3;
  reg [27:0] p21_abs_fraction__2;
  reg [27:0] p21_abs_fraction__3;
  reg [27:0] p21_abs_fraction__4;
  reg [27:0] p21_abs_fraction__5;
  reg p21_ne_9428;
  reg p21_ne_9429;
  reg p21_ne_9430;
  reg p21_ne_9431;
  reg p21_nor_9242;
  reg p21_nor_9245;
  reg p21_is_result_nan__7;
  reg p21_is_operand_inf__2;
  reg p21_is_result_nan__8;
  reg p21_is_operand_inf__3;
  reg p21_is_result_nan__9;
  reg p21_is_result_nan__10;
  reg p21_result_sign__16;
  reg p21_result_sign__18;
  reg p21_result_sign__21;
  reg p21_result_sign__24;
  always_ff @ (posedge clk) begin
    p21_greater_exp_bexp__2 <= p20_greater_exp_bexp__2;
    p21_greater_exp_bexp__3 <= p20_greater_exp_bexp__3;
    p21_abs_fraction__2 <= p21_abs_fraction__2_comb;
    p21_abs_fraction__3 <= p21_abs_fraction__3_comb;
    p21_abs_fraction__4 <= p21_abs_fraction__4_comb;
    p21_abs_fraction__5 <= p21_abs_fraction__5_comb;
    p21_ne_9428 <= p21_ne_9428_comb;
    p21_ne_9429 <= p21_ne_9429_comb;
    p21_ne_9430 <= p21_ne_9430_comb;
    p21_ne_9431 <= p21_ne_9431_comb;
    p21_nor_9242 <= p20_nor_9242;
    p21_nor_9245 <= p20_nor_9245;
    p21_is_result_nan__7 <= p20_is_result_nan__7;
    p21_is_operand_inf__2 <= p20_is_operand_inf__2;
    p21_is_result_nan__8 <= p20_is_result_nan__8;
    p21_is_operand_inf__3 <= p20_is_operand_inf__3;
    p21_is_result_nan__9 <= p20_is_result_nan__9;
    p21_is_result_nan__10 <= p20_is_result_nan__10;
    p21_result_sign__16 <= p21_result_sign__16_comb;
    p21_result_sign__18 <= p21_result_sign__18_comb;
    p21_result_sign__21 <= p21_result_sign__21_comb;
    p21_result_sign__24 <= p21_result_sign__24_comb;
  end

  // ===== Pipe stage 22:
  wire [27:0] p22_reverse_9508_comb;
  wire [27:0] p22_reverse_9509_comb;
  wire [27:0] p22_reverse_9510_comb;
  wire [27:0] p22_reverse_9511_comb;
  wire [28:0] p22_one_hot_9512_comb;
  wire [28:0] p22_one_hot_9513_comb;
  wire [28:0] p22_one_hot_9514_comb;
  wire [28:0] p22_one_hot_9515_comb;
  wire [4:0] p22_encode_9516_comb;
  wire [4:0] p22_encode_9517_comb;
  wire [4:0] p22_encode_9518_comb;
  wire [4:0] p22_encode_9519_comb;
  wire p22_cancel__2_comb;
  wire p22_cancel__3_comb;
  wire p22_cancel__4_comb;
  wire p22_cancel__5_comb;
  wire p22_result_sign__19_comb;
  wire p22_result_sign__22_comb;
  wire p22_result_sign__25_comb;
  wire p22_result_sign__26_comb;
  assign p22_reverse_9508_comb = {p21_abs_fraction__2[0], p21_abs_fraction__2[1], p21_abs_fraction__2[2], p21_abs_fraction__2[3], p21_abs_fraction__2[4], p21_abs_fraction__2[5], p21_abs_fraction__2[6], p21_abs_fraction__2[7], p21_abs_fraction__2[8], p21_abs_fraction__2[9], p21_abs_fraction__2[10], p21_abs_fraction__2[11], p21_abs_fraction__2[12], p21_abs_fraction__2[13], p21_abs_fraction__2[14], p21_abs_fraction__2[15], p21_abs_fraction__2[16], p21_abs_fraction__2[17], p21_abs_fraction__2[18], p21_abs_fraction__2[19], p21_abs_fraction__2[20], p21_abs_fraction__2[21], p21_abs_fraction__2[22], p21_abs_fraction__2[23], p21_abs_fraction__2[24], p21_abs_fraction__2[25], p21_abs_fraction__2[26], p21_abs_fraction__2[27]};
  assign p22_reverse_9509_comb = {p21_abs_fraction__3[0], p21_abs_fraction__3[1], p21_abs_fraction__3[2], p21_abs_fraction__3[3], p21_abs_fraction__3[4], p21_abs_fraction__3[5], p21_abs_fraction__3[6], p21_abs_fraction__3[7], p21_abs_fraction__3[8], p21_abs_fraction__3[9], p21_abs_fraction__3[10], p21_abs_fraction__3[11], p21_abs_fraction__3[12], p21_abs_fraction__3[13], p21_abs_fraction__3[14], p21_abs_fraction__3[15], p21_abs_fraction__3[16], p21_abs_fraction__3[17], p21_abs_fraction__3[18], p21_abs_fraction__3[19], p21_abs_fraction__3[20], p21_abs_fraction__3[21], p21_abs_fraction__3[22], p21_abs_fraction__3[23], p21_abs_fraction__3[24], p21_abs_fraction__3[25], p21_abs_fraction__3[26], p21_abs_fraction__3[27]};
  assign p22_reverse_9510_comb = {p21_abs_fraction__4[0], p21_abs_fraction__4[1], p21_abs_fraction__4[2], p21_abs_fraction__4[3], p21_abs_fraction__4[4], p21_abs_fraction__4[5], p21_abs_fraction__4[6], p21_abs_fraction__4[7], p21_abs_fraction__4[8], p21_abs_fraction__4[9], p21_abs_fraction__4[10], p21_abs_fraction__4[11], p21_abs_fraction__4[12], p21_abs_fraction__4[13], p21_abs_fraction__4[14], p21_abs_fraction__4[15], p21_abs_fraction__4[16], p21_abs_fraction__4[17], p21_abs_fraction__4[18], p21_abs_fraction__4[19], p21_abs_fraction__4[20], p21_abs_fraction__4[21], p21_abs_fraction__4[22], p21_abs_fraction__4[23], p21_abs_fraction__4[24], p21_abs_fraction__4[25], p21_abs_fraction__4[26], p21_abs_fraction__4[27]};
  assign p22_reverse_9511_comb = {p21_abs_fraction__5[0], p21_abs_fraction__5[1], p21_abs_fraction__5[2], p21_abs_fraction__5[3], p21_abs_fraction__5[4], p21_abs_fraction__5[5], p21_abs_fraction__5[6], p21_abs_fraction__5[7], p21_abs_fraction__5[8], p21_abs_fraction__5[9], p21_abs_fraction__5[10], p21_abs_fraction__5[11], p21_abs_fraction__5[12], p21_abs_fraction__5[13], p21_abs_fraction__5[14], p21_abs_fraction__5[15], p21_abs_fraction__5[16], p21_abs_fraction__5[17], p21_abs_fraction__5[18], p21_abs_fraction__5[19], p21_abs_fraction__5[20], p21_abs_fraction__5[21], p21_abs_fraction__5[22], p21_abs_fraction__5[23], p21_abs_fraction__5[24], p21_abs_fraction__5[25], p21_abs_fraction__5[26], p21_abs_fraction__5[27]};
  assign p22_one_hot_9512_comb = {p22_reverse_9508_comb[27:0] == 28'h000_0000, p22_reverse_9508_comb[27] && p22_reverse_9508_comb[26:0] == 27'h000_0000, p22_reverse_9508_comb[26] && p22_reverse_9508_comb[25:0] == 26'h000_0000, p22_reverse_9508_comb[25] && p22_reverse_9508_comb[24:0] == 25'h000_0000, p22_reverse_9508_comb[24] && p22_reverse_9508_comb[23:0] == 24'h00_0000, p22_reverse_9508_comb[23] && p22_reverse_9508_comb[22:0] == 23'h00_0000, p22_reverse_9508_comb[22] && p22_reverse_9508_comb[21:0] == 22'h00_0000, p22_reverse_9508_comb[21] && p22_reverse_9508_comb[20:0] == 21'h00_0000, p22_reverse_9508_comb[20] && p22_reverse_9508_comb[19:0] == 20'h0_0000, p22_reverse_9508_comb[19] && p22_reverse_9508_comb[18:0] == 19'h0_0000, p22_reverse_9508_comb[18] && p22_reverse_9508_comb[17:0] == 18'h0_0000, p22_reverse_9508_comb[17] && p22_reverse_9508_comb[16:0] == 17'h0_0000, p22_reverse_9508_comb[16] && p22_reverse_9508_comb[15:0] == 16'h0000, p22_reverse_9508_comb[15] && p22_reverse_9508_comb[14:0] == 15'h0000, p22_reverse_9508_comb[14] && p22_reverse_9508_comb[13:0] == 14'h0000, p22_reverse_9508_comb[13] && p22_reverse_9508_comb[12:0] == 13'h0000, p22_reverse_9508_comb[12] && p22_reverse_9508_comb[11:0] == 12'h000, p22_reverse_9508_comb[11] && p22_reverse_9508_comb[10:0] == 11'h000, p22_reverse_9508_comb[10] && p22_reverse_9508_comb[9:0] == 10'h000, p22_reverse_9508_comb[9] && p22_reverse_9508_comb[8:0] == 9'h000, p22_reverse_9508_comb[8] && p22_reverse_9508_comb[7:0] == 8'h00, p22_reverse_9508_comb[7] && p22_reverse_9508_comb[6:0] == 7'h00, p22_reverse_9508_comb[6] && p22_reverse_9508_comb[5:0] == 6'h00, p22_reverse_9508_comb[5] && p22_reverse_9508_comb[4:0] == 5'h00, p22_reverse_9508_comb[4] && p22_reverse_9508_comb[3:0] == 4'h0, p22_reverse_9508_comb[3] && p22_reverse_9508_comb[2:0] == 3'h0, p22_reverse_9508_comb[2] && p22_reverse_9508_comb[1:0] == 2'h0, p22_reverse_9508_comb[1] && !p22_reverse_9508_comb[0], p22_reverse_9508_comb[0]};
  assign p22_one_hot_9513_comb = {p22_reverse_9509_comb[27:0] == 28'h000_0000, p22_reverse_9509_comb[27] && p22_reverse_9509_comb[26:0] == 27'h000_0000, p22_reverse_9509_comb[26] && p22_reverse_9509_comb[25:0] == 26'h000_0000, p22_reverse_9509_comb[25] && p22_reverse_9509_comb[24:0] == 25'h000_0000, p22_reverse_9509_comb[24] && p22_reverse_9509_comb[23:0] == 24'h00_0000, p22_reverse_9509_comb[23] && p22_reverse_9509_comb[22:0] == 23'h00_0000, p22_reverse_9509_comb[22] && p22_reverse_9509_comb[21:0] == 22'h00_0000, p22_reverse_9509_comb[21] && p22_reverse_9509_comb[20:0] == 21'h00_0000, p22_reverse_9509_comb[20] && p22_reverse_9509_comb[19:0] == 20'h0_0000, p22_reverse_9509_comb[19] && p22_reverse_9509_comb[18:0] == 19'h0_0000, p22_reverse_9509_comb[18] && p22_reverse_9509_comb[17:0] == 18'h0_0000, p22_reverse_9509_comb[17] && p22_reverse_9509_comb[16:0] == 17'h0_0000, p22_reverse_9509_comb[16] && p22_reverse_9509_comb[15:0] == 16'h0000, p22_reverse_9509_comb[15] && p22_reverse_9509_comb[14:0] == 15'h0000, p22_reverse_9509_comb[14] && p22_reverse_9509_comb[13:0] == 14'h0000, p22_reverse_9509_comb[13] && p22_reverse_9509_comb[12:0] == 13'h0000, p22_reverse_9509_comb[12] && p22_reverse_9509_comb[11:0] == 12'h000, p22_reverse_9509_comb[11] && p22_reverse_9509_comb[10:0] == 11'h000, p22_reverse_9509_comb[10] && p22_reverse_9509_comb[9:0] == 10'h000, p22_reverse_9509_comb[9] && p22_reverse_9509_comb[8:0] == 9'h000, p22_reverse_9509_comb[8] && p22_reverse_9509_comb[7:0] == 8'h00, p22_reverse_9509_comb[7] && p22_reverse_9509_comb[6:0] == 7'h00, p22_reverse_9509_comb[6] && p22_reverse_9509_comb[5:0] == 6'h00, p22_reverse_9509_comb[5] && p22_reverse_9509_comb[4:0] == 5'h00, p22_reverse_9509_comb[4] && p22_reverse_9509_comb[3:0] == 4'h0, p22_reverse_9509_comb[3] && p22_reverse_9509_comb[2:0] == 3'h0, p22_reverse_9509_comb[2] && p22_reverse_9509_comb[1:0] == 2'h0, p22_reverse_9509_comb[1] && !p22_reverse_9509_comb[0], p22_reverse_9509_comb[0]};
  assign p22_one_hot_9514_comb = {p22_reverse_9510_comb[27:0] == 28'h000_0000, p22_reverse_9510_comb[27] && p22_reverse_9510_comb[26:0] == 27'h000_0000, p22_reverse_9510_comb[26] && p22_reverse_9510_comb[25:0] == 26'h000_0000, p22_reverse_9510_comb[25] && p22_reverse_9510_comb[24:0] == 25'h000_0000, p22_reverse_9510_comb[24] && p22_reverse_9510_comb[23:0] == 24'h00_0000, p22_reverse_9510_comb[23] && p22_reverse_9510_comb[22:0] == 23'h00_0000, p22_reverse_9510_comb[22] && p22_reverse_9510_comb[21:0] == 22'h00_0000, p22_reverse_9510_comb[21] && p22_reverse_9510_comb[20:0] == 21'h00_0000, p22_reverse_9510_comb[20] && p22_reverse_9510_comb[19:0] == 20'h0_0000, p22_reverse_9510_comb[19] && p22_reverse_9510_comb[18:0] == 19'h0_0000, p22_reverse_9510_comb[18] && p22_reverse_9510_comb[17:0] == 18'h0_0000, p22_reverse_9510_comb[17] && p22_reverse_9510_comb[16:0] == 17'h0_0000, p22_reverse_9510_comb[16] && p22_reverse_9510_comb[15:0] == 16'h0000, p22_reverse_9510_comb[15] && p22_reverse_9510_comb[14:0] == 15'h0000, p22_reverse_9510_comb[14] && p22_reverse_9510_comb[13:0] == 14'h0000, p22_reverse_9510_comb[13] && p22_reverse_9510_comb[12:0] == 13'h0000, p22_reverse_9510_comb[12] && p22_reverse_9510_comb[11:0] == 12'h000, p22_reverse_9510_comb[11] && p22_reverse_9510_comb[10:0] == 11'h000, p22_reverse_9510_comb[10] && p22_reverse_9510_comb[9:0] == 10'h000, p22_reverse_9510_comb[9] && p22_reverse_9510_comb[8:0] == 9'h000, p22_reverse_9510_comb[8] && p22_reverse_9510_comb[7:0] == 8'h00, p22_reverse_9510_comb[7] && p22_reverse_9510_comb[6:0] == 7'h00, p22_reverse_9510_comb[6] && p22_reverse_9510_comb[5:0] == 6'h00, p22_reverse_9510_comb[5] && p22_reverse_9510_comb[4:0] == 5'h00, p22_reverse_9510_comb[4] && p22_reverse_9510_comb[3:0] == 4'h0, p22_reverse_9510_comb[3] && p22_reverse_9510_comb[2:0] == 3'h0, p22_reverse_9510_comb[2] && p22_reverse_9510_comb[1:0] == 2'h0, p22_reverse_9510_comb[1] && !p22_reverse_9510_comb[0], p22_reverse_9510_comb[0]};
  assign p22_one_hot_9515_comb = {p22_reverse_9511_comb[27:0] == 28'h000_0000, p22_reverse_9511_comb[27] && p22_reverse_9511_comb[26:0] == 27'h000_0000, p22_reverse_9511_comb[26] && p22_reverse_9511_comb[25:0] == 26'h000_0000, p22_reverse_9511_comb[25] && p22_reverse_9511_comb[24:0] == 25'h000_0000, p22_reverse_9511_comb[24] && p22_reverse_9511_comb[23:0] == 24'h00_0000, p22_reverse_9511_comb[23] && p22_reverse_9511_comb[22:0] == 23'h00_0000, p22_reverse_9511_comb[22] && p22_reverse_9511_comb[21:0] == 22'h00_0000, p22_reverse_9511_comb[21] && p22_reverse_9511_comb[20:0] == 21'h00_0000, p22_reverse_9511_comb[20] && p22_reverse_9511_comb[19:0] == 20'h0_0000, p22_reverse_9511_comb[19] && p22_reverse_9511_comb[18:0] == 19'h0_0000, p22_reverse_9511_comb[18] && p22_reverse_9511_comb[17:0] == 18'h0_0000, p22_reverse_9511_comb[17] && p22_reverse_9511_comb[16:0] == 17'h0_0000, p22_reverse_9511_comb[16] && p22_reverse_9511_comb[15:0] == 16'h0000, p22_reverse_9511_comb[15] && p22_reverse_9511_comb[14:0] == 15'h0000, p22_reverse_9511_comb[14] && p22_reverse_9511_comb[13:0] == 14'h0000, p22_reverse_9511_comb[13] && p22_reverse_9511_comb[12:0] == 13'h0000, p22_reverse_9511_comb[12] && p22_reverse_9511_comb[11:0] == 12'h000, p22_reverse_9511_comb[11] && p22_reverse_9511_comb[10:0] == 11'h000, p22_reverse_9511_comb[10] && p22_reverse_9511_comb[9:0] == 10'h000, p22_reverse_9511_comb[9] && p22_reverse_9511_comb[8:0] == 9'h000, p22_reverse_9511_comb[8] && p22_reverse_9511_comb[7:0] == 8'h00, p22_reverse_9511_comb[7] && p22_reverse_9511_comb[6:0] == 7'h00, p22_reverse_9511_comb[6] && p22_reverse_9511_comb[5:0] == 6'h00, p22_reverse_9511_comb[5] && p22_reverse_9511_comb[4:0] == 5'h00, p22_reverse_9511_comb[4] && p22_reverse_9511_comb[3:0] == 4'h0, p22_reverse_9511_comb[3] && p22_reverse_9511_comb[2:0] == 3'h0, p22_reverse_9511_comb[2] && p22_reverse_9511_comb[1:0] == 2'h0, p22_reverse_9511_comb[1] && !p22_reverse_9511_comb[0], p22_reverse_9511_comb[0]};
  assign p22_encode_9516_comb = {p22_one_hot_9512_comb[16] | p22_one_hot_9512_comb[17] | p22_one_hot_9512_comb[18] | p22_one_hot_9512_comb[19] | p22_one_hot_9512_comb[20] | p22_one_hot_9512_comb[21] | p22_one_hot_9512_comb[22] | p22_one_hot_9512_comb[23] | p22_one_hot_9512_comb[24] | p22_one_hot_9512_comb[25] | p22_one_hot_9512_comb[26] | p22_one_hot_9512_comb[27] | p22_one_hot_9512_comb[28], p22_one_hot_9512_comb[8] | p22_one_hot_9512_comb[9] | p22_one_hot_9512_comb[10] | p22_one_hot_9512_comb[11] | p22_one_hot_9512_comb[12] | p22_one_hot_9512_comb[13] | p22_one_hot_9512_comb[14] | p22_one_hot_9512_comb[15] | p22_one_hot_9512_comb[24] | p22_one_hot_9512_comb[25] | p22_one_hot_9512_comb[26] | p22_one_hot_9512_comb[27] | p22_one_hot_9512_comb[28], p22_one_hot_9512_comb[4] | p22_one_hot_9512_comb[5] | p22_one_hot_9512_comb[6] | p22_one_hot_9512_comb[7] | p22_one_hot_9512_comb[12] | p22_one_hot_9512_comb[13] | p22_one_hot_9512_comb[14] | p22_one_hot_9512_comb[15] | p22_one_hot_9512_comb[20] | p22_one_hot_9512_comb[21] | p22_one_hot_9512_comb[22] | p22_one_hot_9512_comb[23] | p22_one_hot_9512_comb[28], p22_one_hot_9512_comb[2] | p22_one_hot_9512_comb[3] | p22_one_hot_9512_comb[6] | p22_one_hot_9512_comb[7] | p22_one_hot_9512_comb[10] | p22_one_hot_9512_comb[11] | p22_one_hot_9512_comb[14] | p22_one_hot_9512_comb[15] | p22_one_hot_9512_comb[18] | p22_one_hot_9512_comb[19] | p22_one_hot_9512_comb[22] | p22_one_hot_9512_comb[23] | p22_one_hot_9512_comb[26] | p22_one_hot_9512_comb[27], p22_one_hot_9512_comb[1] | p22_one_hot_9512_comb[3] | p22_one_hot_9512_comb[5] | p22_one_hot_9512_comb[7] | p22_one_hot_9512_comb[9] | p22_one_hot_9512_comb[11] | p22_one_hot_9512_comb[13] | p22_one_hot_9512_comb[15] | p22_one_hot_9512_comb[17] | p22_one_hot_9512_comb[19] | p22_one_hot_9512_comb[21] | p22_one_hot_9512_comb[23] | p22_one_hot_9512_comb[25] | p22_one_hot_9512_comb[27]};
  assign p22_encode_9517_comb = {p22_one_hot_9513_comb[16] | p22_one_hot_9513_comb[17] | p22_one_hot_9513_comb[18] | p22_one_hot_9513_comb[19] | p22_one_hot_9513_comb[20] | p22_one_hot_9513_comb[21] | p22_one_hot_9513_comb[22] | p22_one_hot_9513_comb[23] | p22_one_hot_9513_comb[24] | p22_one_hot_9513_comb[25] | p22_one_hot_9513_comb[26] | p22_one_hot_9513_comb[27] | p22_one_hot_9513_comb[28], p22_one_hot_9513_comb[8] | p22_one_hot_9513_comb[9] | p22_one_hot_9513_comb[10] | p22_one_hot_9513_comb[11] | p22_one_hot_9513_comb[12] | p22_one_hot_9513_comb[13] | p22_one_hot_9513_comb[14] | p22_one_hot_9513_comb[15] | p22_one_hot_9513_comb[24] | p22_one_hot_9513_comb[25] | p22_one_hot_9513_comb[26] | p22_one_hot_9513_comb[27] | p22_one_hot_9513_comb[28], p22_one_hot_9513_comb[4] | p22_one_hot_9513_comb[5] | p22_one_hot_9513_comb[6] | p22_one_hot_9513_comb[7] | p22_one_hot_9513_comb[12] | p22_one_hot_9513_comb[13] | p22_one_hot_9513_comb[14] | p22_one_hot_9513_comb[15] | p22_one_hot_9513_comb[20] | p22_one_hot_9513_comb[21] | p22_one_hot_9513_comb[22] | p22_one_hot_9513_comb[23] | p22_one_hot_9513_comb[28], p22_one_hot_9513_comb[2] | p22_one_hot_9513_comb[3] | p22_one_hot_9513_comb[6] | p22_one_hot_9513_comb[7] | p22_one_hot_9513_comb[10] | p22_one_hot_9513_comb[11] | p22_one_hot_9513_comb[14] | p22_one_hot_9513_comb[15] | p22_one_hot_9513_comb[18] | p22_one_hot_9513_comb[19] | p22_one_hot_9513_comb[22] | p22_one_hot_9513_comb[23] | p22_one_hot_9513_comb[26] | p22_one_hot_9513_comb[27], p22_one_hot_9513_comb[1] | p22_one_hot_9513_comb[3] | p22_one_hot_9513_comb[5] | p22_one_hot_9513_comb[7] | p22_one_hot_9513_comb[9] | p22_one_hot_9513_comb[11] | p22_one_hot_9513_comb[13] | p22_one_hot_9513_comb[15] | p22_one_hot_9513_comb[17] | p22_one_hot_9513_comb[19] | p22_one_hot_9513_comb[21] | p22_one_hot_9513_comb[23] | p22_one_hot_9513_comb[25] | p22_one_hot_9513_comb[27]};
  assign p22_encode_9518_comb = {p22_one_hot_9514_comb[16] | p22_one_hot_9514_comb[17] | p22_one_hot_9514_comb[18] | p22_one_hot_9514_comb[19] | p22_one_hot_9514_comb[20] | p22_one_hot_9514_comb[21] | p22_one_hot_9514_comb[22] | p22_one_hot_9514_comb[23] | p22_one_hot_9514_comb[24] | p22_one_hot_9514_comb[25] | p22_one_hot_9514_comb[26] | p22_one_hot_9514_comb[27] | p22_one_hot_9514_comb[28], p22_one_hot_9514_comb[8] | p22_one_hot_9514_comb[9] | p22_one_hot_9514_comb[10] | p22_one_hot_9514_comb[11] | p22_one_hot_9514_comb[12] | p22_one_hot_9514_comb[13] | p22_one_hot_9514_comb[14] | p22_one_hot_9514_comb[15] | p22_one_hot_9514_comb[24] | p22_one_hot_9514_comb[25] | p22_one_hot_9514_comb[26] | p22_one_hot_9514_comb[27] | p22_one_hot_9514_comb[28], p22_one_hot_9514_comb[4] | p22_one_hot_9514_comb[5] | p22_one_hot_9514_comb[6] | p22_one_hot_9514_comb[7] | p22_one_hot_9514_comb[12] | p22_one_hot_9514_comb[13] | p22_one_hot_9514_comb[14] | p22_one_hot_9514_comb[15] | p22_one_hot_9514_comb[20] | p22_one_hot_9514_comb[21] | p22_one_hot_9514_comb[22] | p22_one_hot_9514_comb[23] | p22_one_hot_9514_comb[28], p22_one_hot_9514_comb[2] | p22_one_hot_9514_comb[3] | p22_one_hot_9514_comb[6] | p22_one_hot_9514_comb[7] | p22_one_hot_9514_comb[10] | p22_one_hot_9514_comb[11] | p22_one_hot_9514_comb[14] | p22_one_hot_9514_comb[15] | p22_one_hot_9514_comb[18] | p22_one_hot_9514_comb[19] | p22_one_hot_9514_comb[22] | p22_one_hot_9514_comb[23] | p22_one_hot_9514_comb[26] | p22_one_hot_9514_comb[27], p22_one_hot_9514_comb[1] | p22_one_hot_9514_comb[3] | p22_one_hot_9514_comb[5] | p22_one_hot_9514_comb[7] | p22_one_hot_9514_comb[9] | p22_one_hot_9514_comb[11] | p22_one_hot_9514_comb[13] | p22_one_hot_9514_comb[15] | p22_one_hot_9514_comb[17] | p22_one_hot_9514_comb[19] | p22_one_hot_9514_comb[21] | p22_one_hot_9514_comb[23] | p22_one_hot_9514_comb[25] | p22_one_hot_9514_comb[27]};
  assign p22_encode_9519_comb = {p22_one_hot_9515_comb[16] | p22_one_hot_9515_comb[17] | p22_one_hot_9515_comb[18] | p22_one_hot_9515_comb[19] | p22_one_hot_9515_comb[20] | p22_one_hot_9515_comb[21] | p22_one_hot_9515_comb[22] | p22_one_hot_9515_comb[23] | p22_one_hot_9515_comb[24] | p22_one_hot_9515_comb[25] | p22_one_hot_9515_comb[26] | p22_one_hot_9515_comb[27] | p22_one_hot_9515_comb[28], p22_one_hot_9515_comb[8] | p22_one_hot_9515_comb[9] | p22_one_hot_9515_comb[10] | p22_one_hot_9515_comb[11] | p22_one_hot_9515_comb[12] | p22_one_hot_9515_comb[13] | p22_one_hot_9515_comb[14] | p22_one_hot_9515_comb[15] | p22_one_hot_9515_comb[24] | p22_one_hot_9515_comb[25] | p22_one_hot_9515_comb[26] | p22_one_hot_9515_comb[27] | p22_one_hot_9515_comb[28], p22_one_hot_9515_comb[4] | p22_one_hot_9515_comb[5] | p22_one_hot_9515_comb[6] | p22_one_hot_9515_comb[7] | p22_one_hot_9515_comb[12] | p22_one_hot_9515_comb[13] | p22_one_hot_9515_comb[14] | p22_one_hot_9515_comb[15] | p22_one_hot_9515_comb[20] | p22_one_hot_9515_comb[21] | p22_one_hot_9515_comb[22] | p22_one_hot_9515_comb[23] | p22_one_hot_9515_comb[28], p22_one_hot_9515_comb[2] | p22_one_hot_9515_comb[3] | p22_one_hot_9515_comb[6] | p22_one_hot_9515_comb[7] | p22_one_hot_9515_comb[10] | p22_one_hot_9515_comb[11] | p22_one_hot_9515_comb[14] | p22_one_hot_9515_comb[15] | p22_one_hot_9515_comb[18] | p22_one_hot_9515_comb[19] | p22_one_hot_9515_comb[22] | p22_one_hot_9515_comb[23] | p22_one_hot_9515_comb[26] | p22_one_hot_9515_comb[27], p22_one_hot_9515_comb[1] | p22_one_hot_9515_comb[3] | p22_one_hot_9515_comb[5] | p22_one_hot_9515_comb[7] | p22_one_hot_9515_comb[9] | p22_one_hot_9515_comb[11] | p22_one_hot_9515_comb[13] | p22_one_hot_9515_comb[15] | p22_one_hot_9515_comb[17] | p22_one_hot_9515_comb[19] | p22_one_hot_9515_comb[21] | p22_one_hot_9515_comb[23] | p22_one_hot_9515_comb[25] | p22_one_hot_9515_comb[27]};
  assign p22_cancel__2_comb = p22_encode_9516_comb[1] | p22_encode_9516_comb[2] | p22_encode_9516_comb[3] | p22_encode_9516_comb[4];
  assign p22_cancel__3_comb = p22_encode_9517_comb[1] | p22_encode_9517_comb[2] | p22_encode_9517_comb[3] | p22_encode_9517_comb[4];
  assign p22_cancel__4_comb = p22_encode_9518_comb[1] | p22_encode_9518_comb[2] | p22_encode_9518_comb[3] | p22_encode_9518_comb[4];
  assign p22_cancel__5_comb = p22_encode_9519_comb[1] | p22_encode_9519_comb[2] | p22_encode_9519_comb[3] | p22_encode_9519_comb[4];
  assign p22_result_sign__19_comb = ~p21_is_result_nan__7 & p21_result_sign__16;
  assign p22_result_sign__22_comb = ~p21_is_result_nan__8 & p21_result_sign__18;
  assign p22_result_sign__25_comb = ~p21_is_result_nan__9 & p21_result_sign__21;
  assign p22_result_sign__26_comb = ~p21_is_result_nan__10 & p21_result_sign__24;

  // Registers for pipe stage 22:
  reg [7:0] p22_greater_exp_bexp__2;
  reg [7:0] p22_greater_exp_bexp__3;
  reg [27:0] p22_abs_fraction__2;
  reg [27:0] p22_abs_fraction__3;
  reg [27:0] p22_abs_fraction__4;
  reg [27:0] p22_abs_fraction__5;
  reg [4:0] p22_encode_9516;
  reg [4:0] p22_encode_9517;
  reg [4:0] p22_encode_9518;
  reg [4:0] p22_encode_9519;
  reg p22_cancel__2;
  reg p22_cancel__3;
  reg p22_cancel__4;
  reg p22_cancel__5;
  reg p22_ne_9428;
  reg p22_ne_9429;
  reg p22_ne_9430;
  reg p22_ne_9431;
  reg p22_nor_9242;
  reg p22_nor_9245;
  reg p22_is_result_nan__7;
  reg p22_is_operand_inf__2;
  reg p22_is_result_nan__8;
  reg p22_is_operand_inf__3;
  reg p22_is_result_nan__9;
  reg p22_is_result_nan__10;
  reg p22_result_sign__19;
  reg p22_result_sign__22;
  reg p22_result_sign__25;
  reg p22_result_sign__26;
  always_ff @ (posedge clk) begin
    p22_greater_exp_bexp__2 <= p21_greater_exp_bexp__2;
    p22_greater_exp_bexp__3 <= p21_greater_exp_bexp__3;
    p22_abs_fraction__2 <= p21_abs_fraction__2;
    p22_abs_fraction__3 <= p21_abs_fraction__3;
    p22_abs_fraction__4 <= p21_abs_fraction__4;
    p22_abs_fraction__5 <= p21_abs_fraction__5;
    p22_encode_9516 <= p22_encode_9516_comb;
    p22_encode_9517 <= p22_encode_9517_comb;
    p22_encode_9518 <= p22_encode_9518_comb;
    p22_encode_9519 <= p22_encode_9519_comb;
    p22_cancel__2 <= p22_cancel__2_comb;
    p22_cancel__3 <= p22_cancel__3_comb;
    p22_cancel__4 <= p22_cancel__4_comb;
    p22_cancel__5 <= p22_cancel__5_comb;
    p22_ne_9428 <= p21_ne_9428;
    p22_ne_9429 <= p21_ne_9429;
    p22_ne_9430 <= p21_ne_9430;
    p22_ne_9431 <= p21_ne_9431;
    p22_nor_9242 <= p21_nor_9242;
    p22_nor_9245 <= p21_nor_9245;
    p22_is_result_nan__7 <= p21_is_result_nan__7;
    p22_is_operand_inf__2 <= p21_is_operand_inf__2;
    p22_is_result_nan__8 <= p21_is_result_nan__8;
    p22_is_operand_inf__3 <= p21_is_operand_inf__3;
    p22_is_result_nan__9 <= p21_is_result_nan__9;
    p22_is_result_nan__10 <= p21_is_result_nan__10;
    p22_result_sign__19 <= p22_result_sign__19_comb;
    p22_result_sign__22 <= p22_result_sign__22_comb;
    p22_result_sign__25 <= p22_result_sign__25_comb;
    p22_result_sign__26 <= p22_result_sign__26_comb;
  end

  // ===== Pipe stage 23:
  wire p23_carry_bit__2_comb;
  wire p23_carry_bit__3_comb;
  wire p23_carry_bit__4_comb;
  wire p23_carry_bit__5_comb;
  wire [27:0] p23_leading_zeroes__2_comb;
  wire [27:0] p23_leading_zeroes__3_comb;
  wire [27:0] p23_leading_zeroes__4_comb;
  wire [27:0] p23_leading_zeroes__5_comb;
  wire [26:0] p23_carry_fraction__4_comb;
  wire [27:0] p23_add_9646_comb;
  wire [26:0] p23_carry_fraction__6_comb;
  wire [27:0] p23_add_9653_comb;
  wire [26:0] p23_carry_fraction__8_comb;
  wire [27:0] p23_add_9660_comb;
  wire [26:0] p23_carry_fraction__10_comb;
  wire [27:0] p23_add_9667_comb;
  wire [2:0] p23_concat_9668_comb;
  wire [26:0] p23_carry_fraction__5_comb;
  wire [26:0] p23_cancel_fraction__2_comb;
  wire [2:0] p23_concat_9671_comb;
  wire [26:0] p23_carry_fraction__7_comb;
  wire [26:0] p23_cancel_fraction__3_comb;
  wire [2:0] p23_concat_9674_comb;
  wire [26:0] p23_carry_fraction__9_comb;
  wire [26:0] p23_cancel_fraction__4_comb;
  wire [2:0] p23_concat_9677_comb;
  wire [26:0] p23_carry_fraction__11_comb;
  wire [26:0] p23_cancel_fraction__5_comb;
  wire [26:0] p23_shifted_fraction__2_comb;
  wire [26:0] p23_shifted_fraction__3_comb;
  wire [26:0] p23_shifted_fraction__4_comb;
  wire [26:0] p23_shifted_fraction__5_comb;
  assign p23_carry_bit__2_comb = p22_abs_fraction__2[27];
  assign p23_carry_bit__3_comb = p22_abs_fraction__3[27];
  assign p23_carry_bit__4_comb = p22_abs_fraction__4[27];
  assign p23_carry_bit__5_comb = p22_abs_fraction__5[27];
  assign p23_leading_zeroes__2_comb = {23'h00_0000, p22_encode_9516};
  assign p23_leading_zeroes__3_comb = {23'h00_0000, p22_encode_9517};
  assign p23_leading_zeroes__4_comb = {23'h00_0000, p22_encode_9518};
  assign p23_leading_zeroes__5_comb = {23'h00_0000, p22_encode_9519};
  assign p23_carry_fraction__4_comb = p22_abs_fraction__2[27:1];
  assign p23_add_9646_comb = p23_leading_zeroes__2_comb + 28'hfff_ffff;
  assign p23_carry_fraction__6_comb = p22_abs_fraction__3[27:1];
  assign p23_add_9653_comb = p23_leading_zeroes__3_comb + 28'hfff_ffff;
  assign p23_carry_fraction__8_comb = p22_abs_fraction__4[27:1];
  assign p23_add_9660_comb = p23_leading_zeroes__4_comb + 28'hfff_ffff;
  assign p23_carry_fraction__10_comb = p22_abs_fraction__5[27:1];
  assign p23_add_9667_comb = p23_leading_zeroes__5_comb + 28'hfff_ffff;
  assign p23_concat_9668_comb = {~p23_carry_bit__2_comb & ~p22_cancel__2, ~p23_carry_bit__2_comb & p22_cancel__2, p23_carry_bit__2_comb & ~p22_cancel__2};
  assign p23_carry_fraction__5_comb = p23_carry_fraction__4_comb | {26'h000_0000, p22_abs_fraction__2[0]};
  assign p23_cancel_fraction__2_comb = p23_add_9646_comb >= 28'h000_001b ? 27'h000_0000 : p22_abs_fraction__2[26:0] << p23_add_9646_comb;
  assign p23_concat_9671_comb = {~p23_carry_bit__3_comb & ~p22_cancel__3, ~p23_carry_bit__3_comb & p22_cancel__3, p23_carry_bit__3_comb & ~p22_cancel__3};
  assign p23_carry_fraction__7_comb = p23_carry_fraction__6_comb | {26'h000_0000, p22_abs_fraction__3[0]};
  assign p23_cancel_fraction__3_comb = p23_add_9653_comb >= 28'h000_001b ? 27'h000_0000 : p22_abs_fraction__3[26:0] << p23_add_9653_comb;
  assign p23_concat_9674_comb = {~p23_carry_bit__4_comb & ~p22_cancel__4, ~p23_carry_bit__4_comb & p22_cancel__4, p23_carry_bit__4_comb & ~p22_cancel__4};
  assign p23_carry_fraction__9_comb = p23_carry_fraction__8_comb | {26'h000_0000, p22_abs_fraction__4[0]};
  assign p23_cancel_fraction__4_comb = p23_add_9660_comb >= 28'h000_001b ? 27'h000_0000 : p22_abs_fraction__4[26:0] << p23_add_9660_comb;
  assign p23_concat_9677_comb = {~p23_carry_bit__5_comb & ~p22_cancel__5, ~p23_carry_bit__5_comb & p22_cancel__5, p23_carry_bit__5_comb & ~p22_cancel__5};
  assign p23_carry_fraction__11_comb = p23_carry_fraction__10_comb | {26'h000_0000, p22_abs_fraction__5[0]};
  assign p23_cancel_fraction__5_comb = p23_add_9667_comb >= 28'h000_001b ? 27'h000_0000 : p22_abs_fraction__5[26:0] << p23_add_9667_comb;
  assign p23_shifted_fraction__2_comb = p23_carry_fraction__5_comb & {27{p23_concat_9668_comb[0]}} | p23_cancel_fraction__2_comb & {27{p23_concat_9668_comb[1]}} | p22_abs_fraction__2[26:0] & {27{p23_concat_9668_comb[2]}};
  assign p23_shifted_fraction__3_comb = p23_carry_fraction__7_comb & {27{p23_concat_9671_comb[0]}} | p23_cancel_fraction__3_comb & {27{p23_concat_9671_comb[1]}} | p22_abs_fraction__3[26:0] & {27{p23_concat_9671_comb[2]}};
  assign p23_shifted_fraction__4_comb = p23_carry_fraction__9_comb & {27{p23_concat_9674_comb[0]}} | p23_cancel_fraction__4_comb & {27{p23_concat_9674_comb[1]}} | p22_abs_fraction__4[26:0] & {27{p23_concat_9674_comb[2]}};
  assign p23_shifted_fraction__5_comb = p23_carry_fraction__11_comb & {27{p23_concat_9677_comb[0]}} | p23_cancel_fraction__5_comb & {27{p23_concat_9677_comb[1]}} | p22_abs_fraction__5[26:0] & {27{p23_concat_9677_comb[2]}};

  // Registers for pipe stage 23:
  reg [7:0] p23_greater_exp_bexp__2;
  reg [7:0] p23_greater_exp_bexp__3;
  reg [4:0] p23_encode_9516;
  reg [4:0] p23_encode_9517;
  reg [4:0] p23_encode_9518;
  reg [4:0] p23_encode_9519;
  reg [26:0] p23_shifted_fraction__2;
  reg [26:0] p23_shifted_fraction__3;
  reg [26:0] p23_shifted_fraction__4;
  reg [26:0] p23_shifted_fraction__5;
  reg p23_ne_9428;
  reg p23_ne_9429;
  reg p23_ne_9430;
  reg p23_ne_9431;
  reg p23_nor_9242;
  reg p23_nor_9245;
  reg p23_is_result_nan__7;
  reg p23_is_operand_inf__2;
  reg p23_is_result_nan__8;
  reg p23_is_operand_inf__3;
  reg p23_is_result_nan__9;
  reg p23_is_result_nan__10;
  reg p23_result_sign__19;
  reg p23_result_sign__22;
  reg p23_result_sign__25;
  reg p23_result_sign__26;
  always_ff @ (posedge clk) begin
    p23_greater_exp_bexp__2 <= p22_greater_exp_bexp__2;
    p23_greater_exp_bexp__3 <= p22_greater_exp_bexp__3;
    p23_encode_9516 <= p22_encode_9516;
    p23_encode_9517 <= p22_encode_9517;
    p23_encode_9518 <= p22_encode_9518;
    p23_encode_9519 <= p22_encode_9519;
    p23_shifted_fraction__2 <= p23_shifted_fraction__2_comb;
    p23_shifted_fraction__3 <= p23_shifted_fraction__3_comb;
    p23_shifted_fraction__4 <= p23_shifted_fraction__4_comb;
    p23_shifted_fraction__5 <= p23_shifted_fraction__5_comb;
    p23_ne_9428 <= p22_ne_9428;
    p23_ne_9429 <= p22_ne_9429;
    p23_ne_9430 <= p22_ne_9430;
    p23_ne_9431 <= p22_ne_9431;
    p23_nor_9242 <= p22_nor_9242;
    p23_nor_9245 <= p22_nor_9245;
    p23_is_result_nan__7 <= p22_is_result_nan__7;
    p23_is_operand_inf__2 <= p22_is_operand_inf__2;
    p23_is_result_nan__8 <= p22_is_result_nan__8;
    p23_is_operand_inf__3 <= p22_is_operand_inf__3;
    p23_is_result_nan__9 <= p22_is_result_nan__9;
    p23_is_result_nan__10 <= p22_is_result_nan__10;
    p23_result_sign__19 <= p22_result_sign__19;
    p23_result_sign__22 <= p22_result_sign__22;
    p23_result_sign__25 <= p22_result_sign__25;
    p23_result_sign__26 <= p22_result_sign__26;
  end

  // ===== Pipe stage 24:
  wire [2:0] p24_normal_chunk__2_comb;
  wire [1:0] p24_half_way_chunk__2_comb;
  wire [2:0] p24_normal_chunk__3_comb;
  wire [1:0] p24_half_way_chunk__3_comb;
  wire [2:0] p24_normal_chunk__4_comb;
  wire [1:0] p24_half_way_chunk__4_comb;
  wire [2:0] p24_normal_chunk__5_comb;
  wire [1:0] p24_half_way_chunk__5_comb;
  wire [24:0] p24_add_9771_comb;
  wire [24:0] p24_add_9775_comb;
  wire [24:0] p24_add_9779_comb;
  wire [24:0] p24_add_9783_comb;
  wire p24_do_round_up__7_comb;
  wire p24_do_round_up__8_comb;
  wire p24_do_round_up__9_comb;
  wire p24_do_round_up__10_comb;
  wire [27:0] p24_rounded_fraction__2_comb;
  wire [27:0] p24_rounded_fraction__3_comb;
  wire [27:0] p24_rounded_fraction__4_comb;
  wire [27:0] p24_rounded_fraction__5_comb;
  assign p24_normal_chunk__2_comb = p23_shifted_fraction__2[2:0];
  assign p24_half_way_chunk__2_comb = p23_shifted_fraction__2[3:2];
  assign p24_normal_chunk__3_comb = p23_shifted_fraction__3[2:0];
  assign p24_half_way_chunk__3_comb = p23_shifted_fraction__3[3:2];
  assign p24_normal_chunk__4_comb = p23_shifted_fraction__4[2:0];
  assign p24_half_way_chunk__4_comb = p23_shifted_fraction__4[3:2];
  assign p24_normal_chunk__5_comb = p23_shifted_fraction__5[2:0];
  assign p24_half_way_chunk__5_comb = p23_shifted_fraction__5[3:2];
  assign p24_add_9771_comb = {1'h0, p23_shifted_fraction__2[26:3]} + 25'h000_0001;
  assign p24_add_9775_comb = {1'h0, p23_shifted_fraction__3[26:3]} + 25'h000_0001;
  assign p24_add_9779_comb = {1'h0, p23_shifted_fraction__4[26:3]} + 25'h000_0001;
  assign p24_add_9783_comb = {1'h0, p23_shifted_fraction__5[26:3]} + 25'h000_0001;
  assign p24_do_round_up__7_comb = p24_normal_chunk__2_comb > 3'h4 | p24_half_way_chunk__2_comb == 2'h3;
  assign p24_do_round_up__8_comb = p24_normal_chunk__3_comb > 3'h4 | p24_half_way_chunk__3_comb == 2'h3;
  assign p24_do_round_up__9_comb = p24_normal_chunk__4_comb > 3'h4 | p24_half_way_chunk__4_comb == 2'h3;
  assign p24_do_round_up__10_comb = p24_normal_chunk__5_comb > 3'h4 | p24_half_way_chunk__5_comb == 2'h3;
  assign p24_rounded_fraction__2_comb = p24_do_round_up__7_comb ? {p24_add_9771_comb, p24_normal_chunk__2_comb} : {1'h0, p23_shifted_fraction__2};
  assign p24_rounded_fraction__3_comb = p24_do_round_up__8_comb ? {p24_add_9775_comb, p24_normal_chunk__3_comb} : {1'h0, p23_shifted_fraction__3};
  assign p24_rounded_fraction__4_comb = p24_do_round_up__9_comb ? {p24_add_9779_comb, p24_normal_chunk__4_comb} : {1'h0, p23_shifted_fraction__4};
  assign p24_rounded_fraction__5_comb = p24_do_round_up__10_comb ? {p24_add_9783_comb, p24_normal_chunk__5_comb} : {1'h0, p23_shifted_fraction__5};

  // Registers for pipe stage 24:
  reg [7:0] p24_greater_exp_bexp__2;
  reg [7:0] p24_greater_exp_bexp__3;
  reg [4:0] p24_encode_9516;
  reg [4:0] p24_encode_9517;
  reg [4:0] p24_encode_9518;
  reg [4:0] p24_encode_9519;
  reg [27:0] p24_rounded_fraction__2;
  reg [27:0] p24_rounded_fraction__3;
  reg [27:0] p24_rounded_fraction__4;
  reg [27:0] p24_rounded_fraction__5;
  reg p24_ne_9428;
  reg p24_ne_9429;
  reg p24_ne_9430;
  reg p24_ne_9431;
  reg p24_nor_9242;
  reg p24_nor_9245;
  reg p24_is_result_nan__7;
  reg p24_is_operand_inf__2;
  reg p24_is_result_nan__8;
  reg p24_is_operand_inf__3;
  reg p24_is_result_nan__9;
  reg p24_is_result_nan__10;
  reg p24_result_sign__19;
  reg p24_result_sign__22;
  reg p24_result_sign__25;
  reg p24_result_sign__26;
  always_ff @ (posedge clk) begin
    p24_greater_exp_bexp__2 <= p23_greater_exp_bexp__2;
    p24_greater_exp_bexp__3 <= p23_greater_exp_bexp__3;
    p24_encode_9516 <= p23_encode_9516;
    p24_encode_9517 <= p23_encode_9517;
    p24_encode_9518 <= p23_encode_9518;
    p24_encode_9519 <= p23_encode_9519;
    p24_rounded_fraction__2 <= p24_rounded_fraction__2_comb;
    p24_rounded_fraction__3 <= p24_rounded_fraction__3_comb;
    p24_rounded_fraction__4 <= p24_rounded_fraction__4_comb;
    p24_rounded_fraction__5 <= p24_rounded_fraction__5_comb;
    p24_ne_9428 <= p23_ne_9428;
    p24_ne_9429 <= p23_ne_9429;
    p24_ne_9430 <= p23_ne_9430;
    p24_ne_9431 <= p23_ne_9431;
    p24_nor_9242 <= p23_nor_9242;
    p24_nor_9245 <= p23_nor_9245;
    p24_is_result_nan__7 <= p23_is_result_nan__7;
    p24_is_operand_inf__2 <= p23_is_operand_inf__2;
    p24_is_result_nan__8 <= p23_is_result_nan__8;
    p24_is_operand_inf__3 <= p23_is_operand_inf__3;
    p24_is_result_nan__9 <= p23_is_result_nan__9;
    p24_is_result_nan__10 <= p23_is_result_nan__10;
    p24_result_sign__19 <= p23_result_sign__19;
    p24_result_sign__22 <= p23_result_sign__22;
    p24_result_sign__25 <= p23_result_sign__25;
    p24_result_sign__26 <= p23_result_sign__26;
  end

  // ===== Pipe stage 25:
  wire p25_rounding_carry__2_comb;
  wire p25_rounding_carry__3_comb;
  wire p25_rounding_carry__4_comb;
  wire p25_rounding_carry__5_comb;
  wire [8:0] p25_concat_9862_comb;
  wire [8:0] p25_concat_9864_comb;
  wire [8:0] p25_add_9869_comb;
  wire [8:0] p25_add_9871_comb;
  wire [8:0] p25_add_9873_comb;
  wire [8:0] p25_add_9875_comb;
  wire [2:0] p25_add_9900_comb;
  wire [2:0] p25_add_9901_comb;
  wire [2:0] p25_add_9902_comb;
  wire [2:0] p25_add_9903_comb;
  wire [27:0] p25_shrl_9904_comb;
  wire [27:0] p25_shrl_9905_comb;
  wire [27:0] p25_shrl_9906_comb;
  wire [27:0] p25_shrl_9907_comb;
  wire [9:0] p25_add_9884_comb;
  wire [9:0] p25_add_9885_comb;
  wire [9:0] p25_add_9886_comb;
  wire [9:0] p25_add_9887_comb;
  wire [22:0] p25_result_fraction__19_comb;
  wire [22:0] p25_result_fraction__21_comb;
  wire [22:0] p25_result_fraction__24_comb;
  wire [22:0] p25_result_fraction__27_comb;
  assign p25_rounding_carry__2_comb = p24_rounded_fraction__2[27];
  assign p25_rounding_carry__3_comb = p24_rounded_fraction__3[27];
  assign p25_rounding_carry__4_comb = p24_rounded_fraction__4[27];
  assign p25_rounding_carry__5_comb = p24_rounded_fraction__5[27];
  assign p25_concat_9862_comb = {1'h0, p24_greater_exp_bexp__2};
  assign p25_concat_9864_comb = {1'h0, p24_greater_exp_bexp__3};
  assign p25_add_9869_comb = p25_concat_9862_comb + {8'h00, p25_rounding_carry__2_comb};
  assign p25_add_9871_comb = p25_concat_9864_comb + {8'h00, p25_rounding_carry__3_comb};
  assign p25_add_9873_comb = p25_concat_9862_comb + {8'h00, p25_rounding_carry__4_comb};
  assign p25_add_9875_comb = p25_concat_9864_comb + {8'h00, p25_rounding_carry__5_comb};
  assign p25_add_9900_comb = {2'h0, p25_rounding_carry__2_comb} + 3'h3;
  assign p25_add_9901_comb = {2'h0, p25_rounding_carry__3_comb} + 3'h3;
  assign p25_add_9902_comb = {2'h0, p25_rounding_carry__4_comb} + 3'h3;
  assign p25_add_9903_comb = {2'h0, p25_rounding_carry__5_comb} + 3'h3;
  assign p25_shrl_9904_comb = p24_rounded_fraction__2 >> p25_add_9900_comb;
  assign p25_shrl_9905_comb = p24_rounded_fraction__3 >> p25_add_9901_comb;
  assign p25_shrl_9906_comb = p24_rounded_fraction__4 >> p25_add_9902_comb;
  assign p25_shrl_9907_comb = p24_rounded_fraction__5 >> p25_add_9903_comb;
  assign p25_add_9884_comb = {1'h0, p25_add_9869_comb} + 10'h001;
  assign p25_add_9885_comb = {1'h0, p25_add_9871_comb} + 10'h001;
  assign p25_add_9886_comb = {1'h0, p25_add_9873_comb} + 10'h001;
  assign p25_add_9887_comb = {1'h0, p25_add_9875_comb} + 10'h001;
  assign p25_result_fraction__19_comb = p25_shrl_9904_comb[22:0];
  assign p25_result_fraction__21_comb = p25_shrl_9905_comb[22:0];
  assign p25_result_fraction__24_comb = p25_shrl_9906_comb[22:0];
  assign p25_result_fraction__27_comb = p25_shrl_9907_comb[22:0];

  // Registers for pipe stage 25:
  reg [4:0] p25_encode_9516;
  reg [4:0] p25_encode_9517;
  reg [4:0] p25_encode_9518;
  reg [4:0] p25_encode_9519;
  reg [9:0] p25_add_9884;
  reg p25_ne_9428;
  reg [9:0] p25_add_9885;
  reg p25_ne_9429;
  reg [9:0] p25_add_9886;
  reg p25_ne_9430;
  reg [9:0] p25_add_9887;
  reg p25_ne_9431;
  reg p25_nor_9242;
  reg p25_nor_9245;
  reg p25_is_result_nan__7;
  reg p25_is_operand_inf__2;
  reg [22:0] p25_result_fraction__19;
  reg p25_is_result_nan__8;
  reg p25_is_operand_inf__3;
  reg [22:0] p25_result_fraction__21;
  reg p25_is_result_nan__9;
  reg [22:0] p25_result_fraction__24;
  reg p25_is_result_nan__10;
  reg [22:0] p25_result_fraction__27;
  reg p25_result_sign__19;
  reg p25_result_sign__22;
  reg p25_result_sign__25;
  reg p25_result_sign__26;
  always_ff @ (posedge clk) begin
    p25_encode_9516 <= p24_encode_9516;
    p25_encode_9517 <= p24_encode_9517;
    p25_encode_9518 <= p24_encode_9518;
    p25_encode_9519 <= p24_encode_9519;
    p25_add_9884 <= p25_add_9884_comb;
    p25_ne_9428 <= p24_ne_9428;
    p25_add_9885 <= p25_add_9885_comb;
    p25_ne_9429 <= p24_ne_9429;
    p25_add_9886 <= p25_add_9886_comb;
    p25_ne_9430 <= p24_ne_9430;
    p25_add_9887 <= p25_add_9887_comb;
    p25_ne_9431 <= p24_ne_9431;
    p25_nor_9242 <= p24_nor_9242;
    p25_nor_9245 <= p24_nor_9245;
    p25_is_result_nan__7 <= p24_is_result_nan__7;
    p25_is_operand_inf__2 <= p24_is_operand_inf__2;
    p25_result_fraction__19 <= p25_result_fraction__19_comb;
    p25_is_result_nan__8 <= p24_is_result_nan__8;
    p25_is_operand_inf__3 <= p24_is_operand_inf__3;
    p25_result_fraction__21 <= p25_result_fraction__21_comb;
    p25_is_result_nan__9 <= p24_is_result_nan__9;
    p25_result_fraction__24 <= p25_result_fraction__24_comb;
    p25_is_result_nan__10 <= p24_is_result_nan__10;
    p25_result_fraction__27 <= p25_result_fraction__27_comb;
    p25_result_sign__19 <= p24_result_sign__19;
    p25_result_sign__22 <= p24_result_sign__22;
    p25_result_sign__25 <= p24_result_sign__25;
    p25_result_sign__26 <= p24_result_sign__26;
  end

  // ===== Pipe stage 26:
  wire [9:0] p26_wide_exponent__6_comb;
  wire [9:0] p26_wide_exponent__9_comb;
  wire [9:0] p26_wide_exponent__12_comb;
  wire [9:0] p26_wide_exponent__15_comb;
  wire [9:0] p26_wide_exponent__7_comb;
  wire [9:0] p26_wide_exponent__10_comb;
  wire [9:0] p26_wide_exponent__13_comb;
  wire [9:0] p26_wide_exponent__16_comb;
  wire p26_bit_slice_9988_comb;
  wire p26_bit_slice_9989_comb;
  wire p26_bit_slice_9990_comb;
  wire p26_bit_slice_9991_comb;
  wire [8:0] p26_bit_slice_9992_comb;
  wire [8:0] p26_bit_slice_9993_comb;
  wire [8:0] p26_bit_slice_9994_comb;
  wire [8:0] p26_bit_slice_9995_comb;
  assign p26_wide_exponent__6_comb = p25_add_9884 - {5'h00, p25_encode_9516};
  assign p26_wide_exponent__9_comb = p25_add_9885 - {5'h00, p25_encode_9517};
  assign p26_wide_exponent__12_comb = p25_add_9886 - {5'h00, p25_encode_9518};
  assign p26_wide_exponent__15_comb = p25_add_9887 - {5'h00, p25_encode_9519};
  assign p26_wide_exponent__7_comb = p26_wide_exponent__6_comb & {10{p25_ne_9428}};
  assign p26_wide_exponent__10_comb = p26_wide_exponent__9_comb & {10{p25_ne_9429}};
  assign p26_wide_exponent__13_comb = p26_wide_exponent__12_comb & {10{p25_ne_9430}};
  assign p26_wide_exponent__16_comb = p26_wide_exponent__15_comb & {10{p25_ne_9431}};
  assign p26_bit_slice_9988_comb = p26_wide_exponent__7_comb[9];
  assign p26_bit_slice_9989_comb = p26_wide_exponent__10_comb[9];
  assign p26_bit_slice_9990_comb = p26_wide_exponent__13_comb[9];
  assign p26_bit_slice_9991_comb = p26_wide_exponent__16_comb[9];
  assign p26_bit_slice_9992_comb = p26_wide_exponent__7_comb[8:0];
  assign p26_bit_slice_9993_comb = p26_wide_exponent__10_comb[8:0];
  assign p26_bit_slice_9994_comb = p26_wide_exponent__13_comb[8:0];
  assign p26_bit_slice_9995_comb = p26_wide_exponent__16_comb[8:0];

  // Registers for pipe stage 26:
  reg p26_bit_slice_9988;
  reg p26_bit_slice_9989;
  reg p26_bit_slice_9990;
  reg p26_bit_slice_9991;
  reg [8:0] p26_bit_slice_9992;
  reg [8:0] p26_bit_slice_9993;
  reg [8:0] p26_bit_slice_9994;
  reg [8:0] p26_bit_slice_9995;
  reg p26_nor_9242;
  reg p26_nor_9245;
  reg p26_is_result_nan__7;
  reg p26_is_operand_inf__2;
  reg [22:0] p26_result_fraction__19;
  reg p26_is_result_nan__8;
  reg p26_is_operand_inf__3;
  reg [22:0] p26_result_fraction__21;
  reg p26_is_result_nan__9;
  reg [22:0] p26_result_fraction__24;
  reg p26_is_result_nan__10;
  reg [22:0] p26_result_fraction__27;
  reg p26_result_sign__19;
  reg p26_result_sign__22;
  reg p26_result_sign__25;
  reg p26_result_sign__26;
  always_ff @ (posedge clk) begin
    p26_bit_slice_9988 <= p26_bit_slice_9988_comb;
    p26_bit_slice_9989 <= p26_bit_slice_9989_comb;
    p26_bit_slice_9990 <= p26_bit_slice_9990_comb;
    p26_bit_slice_9991 <= p26_bit_slice_9991_comb;
    p26_bit_slice_9992 <= p26_bit_slice_9992_comb;
    p26_bit_slice_9993 <= p26_bit_slice_9993_comb;
    p26_bit_slice_9994 <= p26_bit_slice_9994_comb;
    p26_bit_slice_9995 <= p26_bit_slice_9995_comb;
    p26_nor_9242 <= p25_nor_9242;
    p26_nor_9245 <= p25_nor_9245;
    p26_is_result_nan__7 <= p25_is_result_nan__7;
    p26_is_operand_inf__2 <= p25_is_operand_inf__2;
    p26_result_fraction__19 <= p25_result_fraction__19;
    p26_is_result_nan__8 <= p25_is_result_nan__8;
    p26_is_operand_inf__3 <= p25_is_operand_inf__3;
    p26_result_fraction__21 <= p25_result_fraction__21;
    p26_is_result_nan__9 <= p25_is_result_nan__9;
    p26_result_fraction__24 <= p25_result_fraction__24;
    p26_is_result_nan__10 <= p25_is_result_nan__10;
    p26_result_fraction__27 <= p25_result_fraction__27;
    p26_result_sign__19 <= p25_result_sign__19;
    p26_result_sign__22 <= p25_result_sign__22;
    p26_result_sign__25 <= p25_result_sign__25;
    p26_result_sign__26 <= p25_result_sign__26;
  end

  // ===== Pipe stage 27:
  wire [8:0] p27_wide_exponent__8_comb;
  wire [8:0] p27_wide_exponent__11_comb;
  wire [8:0] p27_wide_exponent__14_comb;
  wire [8:0] p27_wide_exponent__17_comb;
  wire p27_bit_slice_10063_comb;
  wire p27_bit_slice_10071_comb;
  wire p27_bit_slice_10079_comb;
  wire p27_bit_slice_10087_comb;
  wire p27_bit_slice_10088_comb;
  wire p27_bit_slice_10090_comb;
  wire p27_bit_slice_10092_comb;
  wire p27_bit_slice_10094_comb;
  wire p27_or_10089_comb;
  wire p27_or_10091_comb;
  wire p27_or_10093_comb;
  wire p27_or_10095_comb;
  wire p27_and_10096_comb;
  wire p27_and_10097_comb;
  wire p27_and_10098_comb;
  wire p27_and_10099_comb;
  wire [7:0] p27_bit_slice_10100_comb;
  wire [7:0] p27_bit_slice_10101_comb;
  wire [7:0] p27_bit_slice_10102_comb;
  wire [7:0] p27_bit_slice_10103_comb;
  assign p27_wide_exponent__8_comb = p26_bit_slice_9992 & {9{~p26_bit_slice_9988}};
  assign p27_wide_exponent__11_comb = p26_bit_slice_9993 & {9{~p26_bit_slice_9989}};
  assign p27_wide_exponent__14_comb = p26_bit_slice_9994 & {9{~p26_bit_slice_9990}};
  assign p27_wide_exponent__17_comb = p26_bit_slice_9995 & {9{~p26_bit_slice_9991}};
  assign p27_bit_slice_10063_comb = p27_wide_exponent__8_comb[8];
  assign p27_bit_slice_10071_comb = p27_wide_exponent__11_comb[8];
  assign p27_bit_slice_10079_comb = p27_wide_exponent__14_comb[8];
  assign p27_bit_slice_10087_comb = p27_wide_exponent__17_comb[8];
  assign p27_bit_slice_10088_comb = p27_wide_exponent__8_comb[0];
  assign p27_bit_slice_10090_comb = p27_wide_exponent__11_comb[0];
  assign p27_bit_slice_10092_comb = p27_wide_exponent__14_comb[0];
  assign p27_bit_slice_10094_comb = p27_wide_exponent__17_comb[0];
  assign p27_or_10089_comb = p27_wide_exponent__8_comb[1] | p27_wide_exponent__8_comb[2] | p27_wide_exponent__8_comb[3] | p27_wide_exponent__8_comb[4] | p27_wide_exponent__8_comb[5] | p27_wide_exponent__8_comb[6] | p27_wide_exponent__8_comb[7] | p27_bit_slice_10063_comb;
  assign p27_or_10091_comb = p27_wide_exponent__11_comb[1] | p27_wide_exponent__11_comb[2] | p27_wide_exponent__11_comb[3] | p27_wide_exponent__11_comb[4] | p27_wide_exponent__11_comb[5] | p27_wide_exponent__11_comb[6] | p27_wide_exponent__11_comb[7] | p27_bit_slice_10071_comb;
  assign p27_or_10093_comb = p27_wide_exponent__14_comb[1] | p27_wide_exponent__14_comb[2] | p27_wide_exponent__14_comb[3] | p27_wide_exponent__14_comb[4] | p27_wide_exponent__14_comb[5] | p27_wide_exponent__14_comb[6] | p27_wide_exponent__14_comb[7] | p27_bit_slice_10079_comb;
  assign p27_or_10095_comb = p27_wide_exponent__17_comb[1] | p27_wide_exponent__17_comb[2] | p27_wide_exponent__17_comb[3] | p27_wide_exponent__17_comb[4] | p27_wide_exponent__17_comb[5] | p27_wide_exponent__17_comb[6] | p27_wide_exponent__17_comb[7] | p27_bit_slice_10087_comb;
  assign p27_and_10096_comb = p27_bit_slice_10088_comb & p27_wide_exponent__8_comb[1] & p27_wide_exponent__8_comb[2] & p27_wide_exponent__8_comb[3] & p27_wide_exponent__8_comb[4] & p27_wide_exponent__8_comb[5] & p27_wide_exponent__8_comb[6] & p27_wide_exponent__8_comb[7];
  assign p27_and_10097_comb = p27_bit_slice_10090_comb & p27_wide_exponent__11_comb[1] & p27_wide_exponent__11_comb[2] & p27_wide_exponent__11_comb[3] & p27_wide_exponent__11_comb[4] & p27_wide_exponent__11_comb[5] & p27_wide_exponent__11_comb[6] & p27_wide_exponent__11_comb[7];
  assign p27_and_10098_comb = p27_bit_slice_10092_comb & p27_wide_exponent__14_comb[1] & p27_wide_exponent__14_comb[2] & p27_wide_exponent__14_comb[3] & p27_wide_exponent__14_comb[4] & p27_wide_exponent__14_comb[5] & p27_wide_exponent__14_comb[6] & p27_wide_exponent__14_comb[7];
  assign p27_and_10099_comb = p27_bit_slice_10094_comb & p27_wide_exponent__17_comb[1] & p27_wide_exponent__17_comb[2] & p27_wide_exponent__17_comb[3] & p27_wide_exponent__17_comb[4] & p27_wide_exponent__17_comb[5] & p27_wide_exponent__17_comb[6] & p27_wide_exponent__17_comb[7];
  assign p27_bit_slice_10100_comb = p27_wide_exponent__8_comb[7:0];
  assign p27_bit_slice_10101_comb = p27_wide_exponent__11_comb[7:0];
  assign p27_bit_slice_10102_comb = p27_wide_exponent__14_comb[7:0];
  assign p27_bit_slice_10103_comb = p27_wide_exponent__17_comb[7:0];

  // Registers for pipe stage 27:
  reg p27_bit_slice_10063;
  reg p27_bit_slice_10071;
  reg p27_bit_slice_10079;
  reg p27_bit_slice_10087;
  reg p27_bit_slice_10088;
  reg p27_or_10089;
  reg p27_bit_slice_10090;
  reg p27_or_10091;
  reg p27_bit_slice_10092;
  reg p27_or_10093;
  reg p27_bit_slice_10094;
  reg p27_or_10095;
  reg p27_and_10096;
  reg p27_and_10097;
  reg p27_and_10098;
  reg p27_and_10099;
  reg p27_nor_9242;
  reg p27_nor_9245;
  reg p27_is_result_nan__7;
  reg p27_is_operand_inf__2;
  reg [22:0] p27_result_fraction__19;
  reg p27_is_result_nan__8;
  reg p27_is_operand_inf__3;
  reg [22:0] p27_result_fraction__21;
  reg p27_is_result_nan__9;
  reg [22:0] p27_result_fraction__24;
  reg p27_is_result_nan__10;
  reg [22:0] p27_result_fraction__27;
  reg [7:0] p27_bit_slice_10100;
  reg [7:0] p27_bit_slice_10101;
  reg [7:0] p27_bit_slice_10102;
  reg [7:0] p27_bit_slice_10103;
  reg p27_result_sign__19;
  reg p27_result_sign__22;
  reg p27_result_sign__25;
  reg p27_result_sign__26;
  always_ff @ (posedge clk) begin
    p27_bit_slice_10063 <= p27_bit_slice_10063_comb;
    p27_bit_slice_10071 <= p27_bit_slice_10071_comb;
    p27_bit_slice_10079 <= p27_bit_slice_10079_comb;
    p27_bit_slice_10087 <= p27_bit_slice_10087_comb;
    p27_bit_slice_10088 <= p27_bit_slice_10088_comb;
    p27_or_10089 <= p27_or_10089_comb;
    p27_bit_slice_10090 <= p27_bit_slice_10090_comb;
    p27_or_10091 <= p27_or_10091_comb;
    p27_bit_slice_10092 <= p27_bit_slice_10092_comb;
    p27_or_10093 <= p27_or_10093_comb;
    p27_bit_slice_10094 <= p27_bit_slice_10094_comb;
    p27_or_10095 <= p27_or_10095_comb;
    p27_and_10096 <= p27_and_10096_comb;
    p27_and_10097 <= p27_and_10097_comb;
    p27_and_10098 <= p27_and_10098_comb;
    p27_and_10099 <= p27_and_10099_comb;
    p27_nor_9242 <= p26_nor_9242;
    p27_nor_9245 <= p26_nor_9245;
    p27_is_result_nan__7 <= p26_is_result_nan__7;
    p27_is_operand_inf__2 <= p26_is_operand_inf__2;
    p27_result_fraction__19 <= p26_result_fraction__19;
    p27_is_result_nan__8 <= p26_is_result_nan__8;
    p27_is_operand_inf__3 <= p26_is_operand_inf__3;
    p27_result_fraction__21 <= p26_result_fraction__21;
    p27_is_result_nan__9 <= p26_is_result_nan__9;
    p27_result_fraction__24 <= p26_result_fraction__24;
    p27_is_result_nan__10 <= p26_is_result_nan__10;
    p27_result_fraction__27 <= p26_result_fraction__27;
    p27_bit_slice_10100 <= p27_bit_slice_10100_comb;
    p27_bit_slice_10101 <= p27_bit_slice_10101_comb;
    p27_bit_slice_10102 <= p27_bit_slice_10102_comb;
    p27_bit_slice_10103 <= p27_bit_slice_10103_comb;
    p27_result_sign__19 <= p26_result_sign__19;
    p27_result_sign__22 <= p26_result_sign__22;
    p27_result_sign__25 <= p26_result_sign__25;
    p27_result_sign__26 <= p26_result_sign__26;
  end

  // ===== Pipe stage 28:
  wire p28_nor_10180_comb;
  wire p28_nor_10182_comb;
  wire p28_nor_10184_comb;
  wire p28_nor_10186_comb;
  wire [22:0] p28_sign_ext_10191_comb;
  wire [22:0] p28_sign_ext_10195_comb;
  wire [7:0] p28_high_exp__42_comb;
  wire [22:0] p28_result_fraction__20_comb;
  wire [22:0] p28_nan_fraction__16_comb;
  wire [7:0] p28_high_exp__43_comb;
  wire [22:0] p28_result_fraction__22_comb;
  wire [22:0] p28_nan_fraction__17_comb;
  wire [7:0] p28_high_exp__44_comb;
  wire [22:0] p28_result_fraction__25_comb;
  wire [22:0] p28_nan_fraction__18_comb;
  wire [7:0] p28_high_exp__45_comb;
  wire [22:0] p28_result_fraction__28_comb;
  wire [22:0] p28_nan_fraction__19_comb;
  wire [7:0] p28_result_exponent__3_comb;
  wire [22:0] p28_result_fraction__23_comb;
  wire [7:0] p28_result_exponent__4_comb;
  wire [22:0] p28_result_fraction__26_comb;
  wire [7:0] p28_result_exponent__5_comb;
  wire [22:0] p28_result_fraction__29_comb;
  wire [7:0] p28_result_exponent__6_comb;
  wire [22:0] p28_result_fraction__30_comb;
  assign p28_nor_10180_comb = ~(p27_bit_slice_10063 | p27_and_10096);
  assign p28_nor_10182_comb = ~(p27_bit_slice_10071 | p27_and_10097);
  assign p28_nor_10184_comb = ~(p27_bit_slice_10079 | p27_and_10098);
  assign p28_nor_10186_comb = ~(p27_bit_slice_10087 | p27_and_10099);
  assign p28_sign_ext_10191_comb = {23{p27_nor_9242}};
  assign p28_sign_ext_10195_comb = {23{p27_nor_9245}};
  assign p28_high_exp__42_comb = 8'hff;
  assign p28_result_fraction__20_comb = p27_result_fraction__19 & {23{~(~(p27_or_10089 | p27_bit_slice_10088))}} & {23{p28_nor_10180_comb}} & p28_sign_ext_10191_comb;
  assign p28_nan_fraction__16_comb = 23'h40_0000;
  assign p28_high_exp__43_comb = 8'hff;
  assign p28_result_fraction__22_comb = p27_result_fraction__21 & {23{~(~(p27_or_10091 | p27_bit_slice_10090))}} & {23{p28_nor_10182_comb}} & p28_sign_ext_10195_comb;
  assign p28_nan_fraction__17_comb = 23'h40_0000;
  assign p28_high_exp__44_comb = 8'hff;
  assign p28_result_fraction__25_comb = p27_result_fraction__24 & {23{~(~(p27_or_10093 | p27_bit_slice_10092))}} & {23{p28_nor_10184_comb}} & p28_sign_ext_10191_comb;
  assign p28_nan_fraction__18_comb = 23'h40_0000;
  assign p28_high_exp__45_comb = 8'hff;
  assign p28_result_fraction__28_comb = p27_result_fraction__27 & {23{~(~(p27_or_10095 | p27_bit_slice_10094))}} & {23{p28_nor_10186_comb}} & p28_sign_ext_10195_comb;
  assign p28_nan_fraction__19_comb = 23'h40_0000;
  assign p28_result_exponent__3_comb = p27_is_result_nan__7 | p27_is_operand_inf__2 | ~p28_nor_10180_comb ? p28_high_exp__42_comb : p27_bit_slice_10100;
  assign p28_result_fraction__23_comb = p27_is_result_nan__7 ? p28_nan_fraction__16_comb : p28_result_fraction__20_comb;
  assign p28_result_exponent__4_comb = p27_is_result_nan__8 | p27_is_operand_inf__3 | ~p28_nor_10182_comb ? p28_high_exp__43_comb : p27_bit_slice_10101;
  assign p28_result_fraction__26_comb = p27_is_result_nan__8 ? p28_nan_fraction__17_comb : p28_result_fraction__22_comb;
  assign p28_result_exponent__5_comb = p27_is_result_nan__9 | p27_is_operand_inf__2 | ~p28_nor_10184_comb ? p28_high_exp__44_comb : p27_bit_slice_10102;
  assign p28_result_fraction__29_comb = p27_is_result_nan__9 ? p28_nan_fraction__18_comb : p28_result_fraction__25_comb;
  assign p28_result_exponent__6_comb = p27_is_result_nan__10 | p27_is_operand_inf__3 | ~p28_nor_10186_comb ? p28_high_exp__45_comb : p27_bit_slice_10103;
  assign p28_result_fraction__30_comb = p27_is_result_nan__10 ? p28_nan_fraction__19_comb : p28_result_fraction__28_comb;

  // Registers for pipe stage 28:
  reg p28_result_sign__19;
  reg [7:0] p28_result_exponent__3;
  reg [22:0] p28_result_fraction__23;
  reg p28_result_sign__22;
  reg [7:0] p28_result_exponent__4;
  reg [22:0] p28_result_fraction__26;
  reg p28_result_sign__25;
  reg [7:0] p28_result_exponent__5;
  reg [22:0] p28_result_fraction__29;
  reg p28_result_sign__26;
  reg [7:0] p28_result_exponent__6;
  reg [22:0] p28_result_fraction__30;
  always_ff @ (posedge clk) begin
    p28_result_sign__19 <= p27_result_sign__19;
    p28_result_exponent__3 <= p28_result_exponent__3_comb;
    p28_result_fraction__23 <= p28_result_fraction__23_comb;
    p28_result_sign__22 <= p27_result_sign__22;
    p28_result_exponent__4 <= p28_result_exponent__4_comb;
    p28_result_fraction__26 <= p28_result_fraction__26_comb;
    p28_result_sign__25 <= p27_result_sign__25;
    p28_result_exponent__5 <= p28_result_exponent__5_comb;
    p28_result_fraction__29 <= p28_result_fraction__29_comb;
    p28_result_sign__26 <= p27_result_sign__26;
    p28_result_exponent__6 <= p28_result_exponent__6_comb;
    p28_result_fraction__30 <= p28_result_fraction__30_comb;
  end

  // ===== Pipe stage 29:
  wire [31:0] p29_out0_r_comb;
  wire [31:0] p29_out0_i_comb;
  wire [31:0] p29_out1_r_comb;
  wire [31:0] p29_out1_i_comb;
  wire [127:0] p29_tuple_10254_comb;
  assign p29_out0_r_comb = {p28_result_sign__19, p28_result_exponent__3, p28_result_fraction__23};
  assign p29_out0_i_comb = {p28_result_sign__22, p28_result_exponent__4, p28_result_fraction__26};
  assign p29_out1_r_comb = {p28_result_sign__25, p28_result_exponent__5, p28_result_fraction__29};
  assign p29_out1_i_comb = {p28_result_sign__26, p28_result_exponent__6, p28_result_fraction__30};
  assign p29_tuple_10254_comb = {p29_out0_r_comb, p29_out0_i_comb, p29_out1_r_comb, p29_out1_i_comb};

  // Registers for pipe stage 29:
  reg [127:0] p29_tuple_10254;
  always_ff @ (posedge clk) begin
    p29_tuple_10254 <= p29_tuple_10254_comb;
  end
  assign out = p29_tuple_10254;
endmodule

module Const #(
  parameter WIDTH = 32,
  parameter VALUE = 0
) (
  output wire logic [WIDTH-1:0] out
);
  assign out = VALUE;
endmodule

//// =========== Computation ============

module Add #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] left,
  input wire logic [IN_WIDTH-1:0] right,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = left + right;
endmodule

module Sub #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] left,
  input wire logic [IN_WIDTH-1:0] right,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = left - right;
endmodule

module MultComb #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] left,
  input wire logic [IN_WIDTH-1:0] right,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = left * right;
endmodule

//// =========== Binary Logical Operations ============

module And #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH-1:0] left,
  input wire logic [WIDTH-1:0] right,
  output wire logic [WIDTH-1:0] out
);
  assign out = left & right;
endmodule

module Or #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic [WIDTH-1:0] out
);
  assign out = left | right;
endmodule

module Xor #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic [WIDTH-1:0] out
);
  assign out = left ^ right;
endmodule

module Not #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] in,
  output wire logic [WIDTH-1:0] out
);
  assign out = ~in;
endmodule

//// =========== Comparions ============

module Gt #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left > right;
endmodule

module Eq #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left == right;
endmodule

module Neq #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left != right;
endmodule

module Lt #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left < right;
endmodule

module Gte #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left >= right;
endmodule

module Lte #(
  parameter WIDTH = 32
) (
  input wire logic  [WIDTH-1:0] left,
  input wire logic  [WIDTH-1:0] right,
  output wire logic out
);
  assign out = left <= right;
endmodule

//// =========== Extension ============

module SignExtend #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  parameter EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = {{EXTEND{in[IN_WIDTH-1]}}, in};
endmodule

module ZeroExtend #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  parameter EXTEND = OUT_WIDTH - IN_WIDTH;
  assign out = {{EXTEND{1'b0}}, in};
endmodule

module Extend #(
  parameter IN_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = {OUT_WIDTH{in}};
endmodule

module Concat #(
  parameter LEFT = 32,
  parameter RIGHT = 32,
  parameter OUT = 64
) (
  input wire logic [LEFT-1:0] left,
  input wire logic [RIGHT-1:0] right,
  output wire logic [OUT-1:0] out
);
  assign out = {left, right};
endmodule

//// =========== Select bits ============
module Select #(
  parameter WIDTH = 32,
  parameter POS = 0
) (
  input wire logic [WIDTH-1:0] in,
  output wire logic out
);
  assign out = in[POS];
endmodule

module Slice #(
  parameter IN_WIDTH = 32,
  parameter MSB = 31,
  parameter LSB = 0,
  parameter OUT_WIDTH = 32
) (
  input wire logic [IN_WIDTH-1:0] in,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = in[MSB:LSB];
endmodule

/// =========== Reduction Operations ============
module ReduceAnd #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  output wire logic out
);
  assign out = &in;
endmodule

module ReduceOr #(
  parameter WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  output wire logic out
);
  assign out = |in;
endmodule

/// ========== Shift Operations ============
module ShiftLeft #(
  parameter WIDTH = 32,
  parameter SHIFT_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  input wire logic [SHIFT_WIDTH-1:0] shift,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = in << shift;
endmodule

module ShiftRight #(
  parameter WIDTH = 32,
  parameter SHIFT_WIDTH = 32,
  parameter OUT_WIDTH = 32
) (
  input wire logic [WIDTH-1:0] in,
  input wire logic [SHIFT_WIDTH-1:0] shift,
  output wire logic [OUT_WIDTH-1:0] out
);
  assign out = in >> shift;
endmodule

module ArithShiftRight #(
  parameter WIDTH = 32
) (
  input wire logic signed [WIDTH-1:0] in,
  input wire logic [WIDTH-1:0] shift,
  output wire logic [WIDTH-1:0] out
); 
  assign out = in >>> shift;
endmodule

module Mux #(
  parameter WIDTH = 32
) (
  input wire logic sel,
  input wire logic [WIDTH-1:0] in0,
  input wire logic [WIDTH-1:0] in1,
  output logic [WIDTH-1:0] out
);
  assign out = sel ? in0 : in1;
endmodule
module undef #(
    parameter WIDTH = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = 'x;
endmodule

module std_const #(
    parameter WIDTH = 32,
    parameter VALUE = 32
) (
   output logic [WIDTH-1:0] out
);
assign out = VALUE;
endmodule

module std_wire #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   output logic [WIDTH-1:0] out
);
assign out = in;
endmodule

module std_add #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] left,
   input logic [WIDTH-1:0] right,
   output logic [WIDTH-1:0] out
);
assign out = left + right;
endmodule

module std_reg #(
    parameter WIDTH = 32
) (
   input logic [WIDTH-1:0] in,
   input logic write_en,
   input logic clk,
   input logic reset,
   output logic [WIDTH-1:0] out,
   output logic done
);
always_ff @(posedge clk) begin
    if (reset) begin
       out <= 0;
       done <= 0;
    end else if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else done <= 1'd0;
  end
endmodule

module comp1(
  input logic [31:0] p2,
  output logic [31:0] p3,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp1
wire _guard0 = 1;
assign p3 = p2;
// COMPONENT END: comp1
endmodule
module comp2(
  input logic [63:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp2
logic [63:0] inst0_in;
logic [31:0] inst0_out;
logic [63:0] inst1_in;
logic [31:0] inst1_out;
logic [31:0] inst2_p2;
logic [31:0] inst2_p3;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(64),
    .LSB(32),
    .MSB(63),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(64),
    .LSB(0),
    .MSB(31),
    .OUT_WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp1 inst2 (
    .clk(inst2_clk),
    .p2(inst2_p2),
    .p3(inst2_p3),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p9 = inst0_out;
assign p10 = inst2_p3;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p2 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp2
endmodule
module comp3(
  input logic [95:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp3
logic [95:0] inst0_in;
logic [31:0] inst0_out;
logic [95:0] inst1_in;
logic [63:0] inst1_out;
logic [63:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(96),
    .LSB(64),
    .MSB(95),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(96),
    .LSB(0),
    .MSB(63),
    .OUT_WIDTH(64)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp2 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp3
endmodule
module comp4(
  input logic [127:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp4
logic [127:0] inst0_in;
logic [31:0] inst0_out;
logic [127:0] inst1_in;
logic [95:0] inst1_out;
logic [95:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(128),
    .LSB(96),
    .MSB(127),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(0),
    .MSB(95),
    .OUT_WIDTH(96)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp3 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp4
endmodule
module comp5(
  input logic [159:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp5
logic [159:0] inst0_in;
logic [31:0] inst0_out;
logic [159:0] inst1_in;
logic [127:0] inst1_out;
logic [127:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(160),
    .LSB(128),
    .MSB(159),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(160),
    .LSB(0),
    .MSB(127),
    .OUT_WIDTH(128)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp4 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp5
endmodule
module comp6(
  input logic [191:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp6
logic [191:0] inst0_in;
logic [31:0] inst0_out;
logic [191:0] inst1_in;
logic [159:0] inst1_out;
logic [159:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(192),
    .LSB(160),
    .MSB(191),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(192),
    .LSB(0),
    .MSB(159),
    .OUT_WIDTH(160)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp5 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp6
endmodule
module comp7(
  input logic [223:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp7
logic [223:0] inst0_in;
logic [31:0] inst0_out;
logic [223:0] inst1_in;
logic [191:0] inst1_out;
logic [191:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(224),
    .LSB(192),
    .MSB(223),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(224),
    .LSB(0),
    .MSB(191),
    .OUT_WIDTH(192)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp6 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp7
endmodule
module comp8(
  input logic [255:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp8
logic [255:0] inst0_in;
logic [31:0] inst0_out;
logic [255:0] inst1_in;
logic [223:0] inst1_out;
logic [223:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(256),
    .LSB(224),
    .MSB(255),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(256),
    .LSB(0),
    .MSB(223),
    .OUT_WIDTH(224)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp7 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp8
endmodule
module comp9(
  input logic [287:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp9
logic [287:0] inst0_in;
logic [31:0] inst0_out;
logic [287:0] inst1_in;
logic [255:0] inst1_out;
logic [255:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(288),
    .LSB(256),
    .MSB(287),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(288),
    .LSB(0),
    .MSB(255),
    .OUT_WIDTH(256)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp8 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp9
endmodule
module comp10(
  input logic [319:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp10
logic [319:0] inst0_in;
logic [31:0] inst0_out;
logic [319:0] inst1_in;
logic [287:0] inst1_out;
logic [287:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(320),
    .LSB(288),
    .MSB(319),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(320),
    .LSB(0),
    .MSB(287),
    .OUT_WIDTH(288)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp9 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp10
endmodule
module comp11(
  input logic [351:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp11
logic [351:0] inst0_in;
logic [31:0] inst0_out;
logic [351:0] inst1_in;
logic [319:0] inst1_out;
logic [319:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(352),
    .LSB(320),
    .MSB(351),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(352),
    .LSB(0),
    .MSB(319),
    .OUT_WIDTH(320)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp10 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp11
endmodule
module comp12(
  input logic [383:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp12
logic [383:0] inst0_in;
logic [31:0] inst0_out;
logic [383:0] inst1_in;
logic [351:0] inst1_out;
logic [351:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(384),
    .LSB(352),
    .MSB(383),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(384),
    .LSB(0),
    .MSB(351),
    .OUT_WIDTH(352)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp11 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp12
endmodule
module comp13(
  input logic [415:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp13
logic [415:0] inst0_in;
logic [31:0] inst0_out;
logic [415:0] inst1_in;
logic [383:0] inst1_out;
logic [383:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(416),
    .LSB(384),
    .MSB(415),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(416),
    .LSB(0),
    .MSB(383),
    .OUT_WIDTH(384)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp12 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp13
endmodule
module comp14(
  input logic [447:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp14
logic [447:0] inst0_in;
logic [31:0] inst0_out;
logic [447:0] inst1_in;
logic [415:0] inst1_out;
logic [415:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(448),
    .LSB(416),
    .MSB(447),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(448),
    .LSB(0),
    .MSB(415),
    .OUT_WIDTH(416)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp13 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp14
endmodule
module comp15(
  input logic [479:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp15
logic [479:0] inst0_in;
logic [31:0] inst0_out;
logic [479:0] inst1_in;
logic [447:0] inst1_out;
logic [447:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(480),
    .LSB(448),
    .MSB(479),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(480),
    .LSB(0),
    .MSB(447),
    .OUT_WIDTH(448)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp14 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp15
endmodule
module comp16(
  input logic [511:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp16
logic [511:0] inst0_in;
logic [31:0] inst0_out;
logic [511:0] inst1_in;
logic [479:0] inst1_out;
logic [479:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(512),
    .LSB(480),
    .MSB(511),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(512),
    .LSB(0),
    .MSB(479),
    .OUT_WIDTH(480)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp15 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp16
endmodule
module comp17(
  input logic [543:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp17
logic [543:0] inst0_in;
logic [31:0] inst0_out;
logic [543:0] inst1_in;
logic [511:0] inst1_out;
logic [511:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(544),
    .LSB(512),
    .MSB(543),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(544),
    .LSB(0),
    .MSB(511),
    .OUT_WIDTH(512)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp16 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp17
endmodule
module comp18(
  input logic [575:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp18
logic [575:0] inst0_in;
logic [31:0] inst0_out;
logic [575:0] inst1_in;
logic [543:0] inst1_out;
logic [543:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(576),
    .LSB(544),
    .MSB(575),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(576),
    .LSB(0),
    .MSB(543),
    .OUT_WIDTH(544)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp17 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp18
endmodule
module comp19(
  input logic [607:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp19
logic [607:0] inst0_in;
logic [31:0] inst0_out;
logic [607:0] inst1_in;
logic [575:0] inst1_out;
logic [575:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(608),
    .LSB(576),
    .MSB(607),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(608),
    .LSB(0),
    .MSB(575),
    .OUT_WIDTH(576)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp18 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp19
endmodule
module comp20(
  input logic [639:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp20
logic [639:0] inst0_in;
logic [31:0] inst0_out;
logic [639:0] inst1_in;
logic [607:0] inst1_out;
logic [607:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(640),
    .LSB(608),
    .MSB(639),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(640),
    .LSB(0),
    .MSB(607),
    .OUT_WIDTH(608)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp19 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp20
endmodule
module comp21(
  input logic [671:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp21
logic [671:0] inst0_in;
logic [31:0] inst0_out;
logic [671:0] inst1_in;
logic [639:0] inst1_out;
logic [639:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(672),
    .LSB(640),
    .MSB(671),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(672),
    .LSB(0),
    .MSB(639),
    .OUT_WIDTH(640)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp20 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp21
endmodule
module comp22(
  input logic [703:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp22
logic [703:0] inst0_in;
logic [31:0] inst0_out;
logic [703:0] inst1_in;
logic [671:0] inst1_out;
logic [671:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(704),
    .LSB(672),
    .MSB(703),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(704),
    .LSB(0),
    .MSB(671),
    .OUT_WIDTH(672)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp21 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp22
endmodule
module comp23(
  input logic [735:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp23
logic [735:0] inst0_in;
logic [31:0] inst0_out;
logic [735:0] inst1_in;
logic [703:0] inst1_out;
logic [703:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(736),
    .LSB(704),
    .MSB(735),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(736),
    .LSB(0),
    .MSB(703),
    .OUT_WIDTH(704)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp22 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp23
endmodule
module comp24(
  input logic [767:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp24
logic [767:0] inst0_in;
logic [31:0] inst0_out;
logic [767:0] inst1_in;
logic [735:0] inst1_out;
logic [735:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(768),
    .LSB(736),
    .MSB(767),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(768),
    .LSB(0),
    .MSB(735),
    .OUT_WIDTH(736)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp23 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp24
endmodule
module comp25(
  input logic [799:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp25
logic [799:0] inst0_in;
logic [31:0] inst0_out;
logic [799:0] inst1_in;
logic [767:0] inst1_out;
logic [767:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(800),
    .LSB(768),
    .MSB(799),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(800),
    .LSB(0),
    .MSB(767),
    .OUT_WIDTH(768)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp24 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp25
endmodule
module comp26(
  input logic [831:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp26
logic [831:0] inst0_in;
logic [31:0] inst0_out;
logic [831:0] inst1_in;
logic [799:0] inst1_out;
logic [799:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(832),
    .LSB(800),
    .MSB(831),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(832),
    .LSB(0),
    .MSB(799),
    .OUT_WIDTH(800)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp25 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp26
endmodule
module comp27(
  input logic [863:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp27
logic [863:0] inst0_in;
logic [31:0] inst0_out;
logic [863:0] inst1_in;
logic [831:0] inst1_out;
logic [831:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(864),
    .LSB(832),
    .MSB(863),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(864),
    .LSB(0),
    .MSB(831),
    .OUT_WIDTH(832)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp26 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp27
endmodule
module comp28(
  input logic [895:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp28
logic [895:0] inst0_in;
logic [31:0] inst0_out;
logic [895:0] inst1_in;
logic [863:0] inst1_out;
logic [863:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(896),
    .LSB(864),
    .MSB(895),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(896),
    .LSB(0),
    .MSB(863),
    .OUT_WIDTH(864)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp27 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp28
endmodule
module comp29(
  input logic [927:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp29
logic [927:0] inst0_in;
logic [31:0] inst0_out;
logic [927:0] inst1_in;
logic [895:0] inst1_out;
logic [895:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(928),
    .LSB(896),
    .MSB(927),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(928),
    .LSB(0),
    .MSB(895),
    .OUT_WIDTH(896)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp28 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp29
endmodule
module comp30(
  input logic [959:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp30
logic [959:0] inst0_in;
logic [31:0] inst0_out;
logic [959:0] inst1_in;
logic [927:0] inst1_out;
logic [927:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic inst2_reset;
logic inst2_clk;
Slice # (
    .IN_WIDTH(960),
    .LSB(928),
    .MSB(959),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(960),
    .LSB(0),
    .MSB(927),
    .OUT_WIDTH(928)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp29 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p38 = inst2_p37;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp30
endmodule
module comp31(
  input logic [991:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp31
logic [991:0] inst0_in;
logic [31:0] inst0_out;
logic [991:0] inst1_in;
logic [959:0] inst1_out;
logic [959:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic [31:0] inst2_p38;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(992),
    .LSB(960),
    .MSB(991),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(992),
    .LSB(0),
    .MSB(959),
    .OUT_WIDTH(960)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp30 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p38(inst2_p38),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p38 = inst2_p37;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p39 = inst2_p38;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp31
endmodule
module comp32(
  input logic [1023:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  output logic [31:0] p40,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp32
logic [1023:0] inst0_in;
logic [31:0] inst0_out;
logic [1023:0] inst1_in;
logic [991:0] inst1_out;
logic [991:0] inst2_p8;
logic [31:0] inst2_p9;
logic [31:0] inst2_p10;
logic [31:0] inst2_p11;
logic [31:0] inst2_p12;
logic [31:0] inst2_p13;
logic [31:0] inst2_p14;
logic [31:0] inst2_p15;
logic [31:0] inst2_p16;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic [31:0] inst2_p33;
logic [31:0] inst2_p34;
logic [31:0] inst2_p35;
logic [31:0] inst2_p36;
logic [31:0] inst2_p37;
logic [31:0] inst2_p38;
logic [31:0] inst2_p39;
logic inst2_clk;
logic inst2_reset;
Slice # (
    .IN_WIDTH(1024),
    .LSB(992),
    .MSB(1023),
    .OUT_WIDTH(32)
) inst0 (
    .in(inst0_in),
    .out(inst0_out)
);
Slice # (
    .IN_WIDTH(1024),
    .LSB(0),
    .MSB(991),
    .OUT_WIDTH(992)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
comp31 inst2 (
    .clk(inst2_clk),
    .p10(inst2_p10),
    .p11(inst2_p11),
    .p12(inst2_p12),
    .p13(inst2_p13),
    .p14(inst2_p14),
    .p15(inst2_p15),
    .p16(inst2_p16),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .p33(inst2_p33),
    .p34(inst2_p34),
    .p35(inst2_p35),
    .p36(inst2_p36),
    .p37(inst2_p37),
    .p38(inst2_p38),
    .p39(inst2_p39),
    .p8(inst2_p8),
    .p9(inst2_p9),
    .reset(inst2_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p18;
assign p28 = inst2_p27;
assign p29 = inst2_p28;
assign p38 = inst2_p37;
assign p40 = inst2_p39;
assign p12 = inst2_p11;
assign p16 = inst2_p15;
assign p9 = inst0_out;
assign p15 = inst2_p14;
assign p17 = inst2_p16;
assign p20 = inst2_p19;
assign p21 = inst2_p20;
assign p23 = inst2_p22;
assign p11 = inst2_p10;
assign p25 = inst2_p24;
assign p36 = inst2_p35;
assign p39 = inst2_p38;
assign p10 = inst2_p9;
assign p13 = inst2_p12;
assign p18 = inst2_p17;
assign p30 = inst2_p29;
assign p24 = inst2_p23;
assign p32 = inst2_p31;
assign p14 = inst2_p13;
assign p26 = inst2_p25;
assign p31 = inst2_p30;
assign p27 = inst2_p26;
assign p33 = inst2_p32;
assign p22 = inst2_p21;
assign p34 = inst2_p33;
assign p35 = inst2_p34;
assign p37 = inst2_p36;
assign inst1_in = p8;
assign inst0_in = p8;
assign inst2_clk = clk;
assign inst2_p8 = inst1_out;
assign inst2_reset = reset;
// COMPONENT END: comp32
endmodule
module comp57(
  input logic [1023:0] p4,
  output logic [31:0] p5,
  output logic [31:0] p6,
  output logic [31:0] p7,
  output logic [31:0] p8,
  output logic [31:0] p9,
  output logic [31:0] p10,
  output logic [31:0] p11,
  output logic [31:0] p12,
  output logic [31:0] p13,
  output logic [31:0] p14,
  output logic [31:0] p15,
  output logic [31:0] p16,
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp57
logic [1023:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [31:0] inst0_p38;
logic [31:0] inst0_p39;
logic [31:0] inst0_p40;
logic inst0_clk;
logic inst0_reset;
comp32 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p39(inst0_p39),
    .p40(inst0_p40),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
wire _guard0 = 1;
assign p19 = inst0_p23;
assign p28 = inst0_p32;
assign p29 = inst0_p33;
assign p12 = inst0_p16;
assign p16 = inst0_p20;
assign p6 = inst0_p10;
assign p9 = inst0_p13;
assign p15 = inst0_p19;
assign p17 = inst0_p21;
assign p20 = inst0_p24;
assign p21 = inst0_p25;
assign p23 = inst0_p27;
assign p11 = inst0_p15;
assign p25 = inst0_p29;
assign p36 = inst0_p40;
assign p5 = inst0_p9;
assign p8 = inst0_p12;
assign p10 = inst0_p14;
assign p13 = inst0_p17;
assign p18 = inst0_p22;
assign p30 = inst0_p34;
assign p7 = inst0_p11;
assign p24 = inst0_p28;
assign p32 = inst0_p36;
assign p14 = inst0_p18;
assign p26 = inst0_p30;
assign p31 = inst0_p35;
assign p27 = inst0_p31;
assign p33 = inst0_p37;
assign p22 = inst0_p26;
assign p34 = inst0_p38;
assign p35 = inst0_p39;
assign inst0_clk = clk;
assign inst0_p8 = p4;
assign inst0_reset = reset;
// COMPONENT END: comp57
endmodule
module comp58(
  input logic [31:0] p2,
  output logic [31:0] p3,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp58
wire _guard0 = 1;
assign p3 = p2;
// COMPONENT END: comp58
endmodule
module comp60(
  input logic [31:0] p7,
  input logic [31:0] p8,
  output logic [63:0] p9,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp60
logic [31:0] inst0_p2;
logic [31:0] inst0_p3;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [31:0] inst1_right;
logic [63:0] inst1_out;
comp58 inst0 (
    .clk(inst0_clk),
    .p2(inst0_p2),
    .p3(inst0_p3),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(64),
    .RIGHT(32)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p9 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p3;
assign inst0_clk = clk;
assign inst0_p2 = p8;
assign inst0_reset = reset;
// COMPONENT END: comp60
endmodule
module comp61(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  output logic [95:0] p10,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp61
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [63:0] inst0_p9;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [63:0] inst1_right;
logic [95:0] inst1_out;
comp60 inst0 (
    .clk(inst0_clk),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(96),
    .RIGHT(64)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p10 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p9;
assign inst0_clk = clk;
assign inst0_p8 = p9;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp61
endmodule
module comp62(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  output logic [127:0] p11,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp62
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [95:0] inst0_p10;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [95:0] inst1_right;
logic [127:0] inst1_out;
comp61 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(128),
    .RIGHT(96)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p11 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p10;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p8 = p9;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp62
endmodule
module comp63(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  output logic [159:0] p12,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp63
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [127:0] inst0_p11;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [127:0] inst1_right;
logic [159:0] inst1_out;
comp62 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(160),
    .RIGHT(128)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p12 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p11;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp63
endmodule
module comp64(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  output logic [191:0] p13,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp64
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [159:0] inst0_p12;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [159:0] inst1_right;
logic [191:0] inst1_out;
comp63 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(192),
    .RIGHT(160)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p13 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p12;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp64
endmodule
module comp65(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  output logic [223:0] p14,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp65
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [191:0] inst0_p13;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [191:0] inst1_right;
logic [223:0] inst1_out;
comp64 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(224),
    .RIGHT(192)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p14 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p13;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p7 = p8;
// COMPONENT END: comp65
endmodule
module comp66(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  output logic [255:0] p15,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp66
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [223:0] inst0_p14;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [223:0] inst1_right;
logic [255:0] inst1_out;
comp65 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(256),
    .RIGHT(224)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p15 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p14;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p7 = p8;
// COMPONENT END: comp66
endmodule
module comp67(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  output logic [287:0] p16,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp67
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [255:0] inst0_p15;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [255:0] inst1_right;
logic [287:0] inst1_out;
comp66 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(288),
    .RIGHT(256)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p16 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p15;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp67
endmodule
module comp68(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  output logic [319:0] p17,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp68
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [287:0] inst0_p16;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [287:0] inst1_right;
logic [319:0] inst1_out;
comp67 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(320),
    .RIGHT(288)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p17 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p16;
assign inst0_p12 = p13;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp68
endmodule
module comp69(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [351:0] p18,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp69
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [319:0] inst0_p17;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [319:0] inst1_right;
logic [351:0] inst1_out;
comp68 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(352),
    .RIGHT(320)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p18 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p17;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp69
endmodule
module comp70(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  output logic [383:0] p19,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp70
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [351:0] inst0_p18;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [351:0] inst1_right;
logic [383:0] inst1_out;
comp69 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(384),
    .RIGHT(352)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p19 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p18;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp70
endmodule
module comp71(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  output logic [415:0] p20,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp71
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [383:0] inst0_p19;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [383:0] inst1_right;
logic [415:0] inst1_out;
comp70 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(416),
    .RIGHT(384)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p20 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p19;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp71
endmodule
module comp72(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  output logic [447:0] p21,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp72
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [415:0] inst0_p20;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [415:0] inst1_right;
logic [447:0] inst1_out;
comp71 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(448),
    .RIGHT(416)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p21 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p20;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp72
endmodule
module comp73(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  output logic [479:0] p22,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp73
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [447:0] inst0_p21;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [447:0] inst1_right;
logic [479:0] inst1_out;
comp72 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(480),
    .RIGHT(448)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p22 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p21;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp73
endmodule
module comp74(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  output logic [511:0] p23,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp74
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [479:0] inst0_p22;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [479:0] inst1_right;
logic [511:0] inst1_out;
comp73 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(512),
    .RIGHT(480)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p23 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p22;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
// COMPONENT END: comp74
endmodule
module comp75(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  output logic [543:0] p24,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp75
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [511:0] inst0_p23;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [511:0] inst1_right;
logic [543:0] inst1_out;
comp74 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(544),
    .RIGHT(512)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p24 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p23;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp75
endmodule
module comp76(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  output logic [575:0] p25,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp76
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [543:0] inst0_p24;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [543:0] inst1_right;
logic [575:0] inst1_out;
comp75 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(576),
    .RIGHT(544)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p25 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p24;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp76
endmodule
module comp77(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  output logic [607:0] p26,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp77
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [575:0] inst0_p25;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [575:0] inst1_right;
logic [607:0] inst1_out;
comp76 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(608),
    .RIGHT(576)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p26 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p25;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp77
endmodule
module comp78(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  output logic [639:0] p27,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp78
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [607:0] inst0_p26;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [607:0] inst1_right;
logic [639:0] inst1_out;
comp77 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(640),
    .RIGHT(608)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p27 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p26;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p22 = p23;
// COMPONENT END: comp78
endmodule
module comp79(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  output logic [671:0] p28,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp79
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [639:0] inst0_p27;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [639:0] inst1_right;
logic [671:0] inst1_out;
comp78 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(672),
    .RIGHT(640)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p28 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p27;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p22 = p23;
// COMPONENT END: comp79
endmodule
module comp80(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  output logic [703:0] p29,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp80
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [671:0] inst0_p28;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [671:0] inst1_right;
logic [703:0] inst1_out;
comp79 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(704),
    .RIGHT(672)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p29 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p28;
assign inst0_p19 = p20;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp80
endmodule
module comp81(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  output logic [735:0] p30,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp81
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [703:0] inst0_p29;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [703:0] inst1_right;
logic [735:0] inst1_out;
comp80 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(736),
    .RIGHT(704)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p30 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p29;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp81
endmodule
module comp82(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  output logic [767:0] p31,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp82
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [735:0] inst0_p30;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [735:0] inst1_right;
logic [767:0] inst1_out;
comp81 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(768),
    .RIGHT(736)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p31 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p30;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp82
endmodule
module comp83(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  output logic [799:0] p32,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp83
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [767:0] inst0_p31;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [767:0] inst1_right;
logic [799:0] inst1_out;
comp82 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(800),
    .RIGHT(768)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p32 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p31;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp83
endmodule
module comp39(
  output logic [31:0] p2,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp39
logic [31:0] inst0_out;
Const # (
    .VALUE(621621554),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp39
endmodule
module comp84(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  output logic [831:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp84
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [799:0] inst0_p32;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [799:0] inst1_right;
logic [831:0] inst1_out;
comp83 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(832),
    .RIGHT(800)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p33 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p32;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp84
endmodule
module comp85(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  output logic [863:0] p34,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp85
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [831:0] inst0_p33;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [831:0] inst1_right;
logic [863:0] inst1_out;
comp84 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(864),
    .RIGHT(832)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p34 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p33;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p22 = p23;
// COMPONENT END: comp85
endmodule
module comp86(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  output logic [895:0] p35,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp86
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [863:0] inst0_p34;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [863:0] inst1_right;
logic [895:0] inst1_out;
comp85 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(896),
    .RIGHT(864)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p35 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p34;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
// COMPONENT END: comp86
endmodule
module comp87(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  output logic [927:0] p36,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp87
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [895:0] inst0_p35;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [895:0] inst1_right;
logic [927:0] inst1_out;
comp86 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(928),
    .RIGHT(896)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p36 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p35;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
// COMPONENT END: comp87
endmodule
module comp88(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  output logic [959:0] p37,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp88
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [927:0] inst0_p36;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_left;
logic [927:0] inst1_right;
logic [959:0] inst1_out;
comp87 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(960),
    .RIGHT(928)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p37 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p36;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
assign inst0_p35 = p36;
// COMPONENT END: comp88
endmodule
module comp89(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  input logic [31:0] p37,
  output logic [991:0] p38,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp89
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [959:0] inst0_p37;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [959:0] inst1_right;
logic [991:0] inst1_out;
comp88 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(992),
    .RIGHT(960)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p38 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p37;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p36 = p37;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
assign inst0_p35 = p36;
// COMPONENT END: comp89
endmodule
module comp90(
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  input logic [31:0] p37,
  input logic [31:0] p38,
  output logic [1023:0] p39,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp90
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [991:0] inst0_p38;
logic inst0_reset;
logic inst0_clk;
logic [31:0] inst1_left;
logic [991:0] inst1_right;
logic [1023:0] inst1_out;
comp89 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
Concat # (
    .LEFT(32),
    .OUT(1024),
    .RIGHT(992)
) inst1 (
    .left(inst1_left),
    .out(inst1_out),
    .right(inst1_right)
);
wire _guard0 = 1;
assign p39 = inst1_out;
assign inst1_left = p7;
assign inst1_right = inst0_p38;
assign inst0_p19 = p20;
assign inst0_p28 = p29;
assign inst0_p29 = p30;
assign inst0_p12 = p13;
assign inst0_p16 = p17;
assign inst0_p9 = p10;
assign inst0_p15 = p16;
assign inst0_p17 = p18;
assign inst0_p20 = p21;
assign inst0_p21 = p22;
assign inst0_p23 = p24;
assign inst0_clk = clk;
assign inst0_p11 = p12;
assign inst0_p25 = p26;
assign inst0_p36 = p37;
assign inst0_p8 = p9;
assign inst0_p10 = p11;
assign inst0_reset = reset;
assign inst0_p13 = p14;
assign inst0_p18 = p19;
assign inst0_p30 = p31;
assign inst0_p7 = p8;
assign inst0_p24 = p25;
assign inst0_p32 = p33;
assign inst0_p14 = p15;
assign inst0_p26 = p27;
assign inst0_p31 = p32;
assign inst0_p27 = p28;
assign inst0_p33 = p34;
assign inst0_p22 = p23;
assign inst0_p34 = p35;
assign inst0_p35 = p36;
assign inst0_p37 = p38;
// COMPONENT END: comp90
endmodule
module comp46(
  output logic [31:0] p4,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp46
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1083407522),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp46
endmodule
module comp42(
  output logic [31:0] p4,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp42
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1094455531),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp42
endmodule
module comp44(
  output logic [31:0] p4,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp44
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1087044365),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp44
endmodule
module comp43(
  output logic [31:0] p2,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp43
logic [31:0] inst0_out;
Const # (
    .VALUE(1060439283),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp43
endmodule
module comp40(
  output logic [31:0] p2,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp40
logic [31:0] inst0_out;
Const # (
    .VALUE(1064076126),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp40
endmodule
module comp38(
  output logic [31:0] p2,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp38
logic [31:0] inst0_out;
Const # (
    .VALUE(1065353216),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp38
endmodule
module comp45(
  output logic [31:0] p2,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp45
logic [31:0] inst0_out;
Const # (
    .VALUE(1053028117),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp45
endmodule
module comp48(
  output logic [31:0] p4,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp48
logic [31:0] inst0_out;
logic [31:0] inst1_in;
logic [31:0] inst1_out;
Const # (
    .VALUE(1082130432),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
Neg # (
    .WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
wire _guard0 = 1;
assign p4 = inst1_out;
assign inst1_in = inst0_out;
// COMPONENT END: comp48
endmodule
module comp47(
  output logic [31:0] p2,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp47
logic [31:0] inst0_out;
Const # (
    .VALUE(613232946),
    .WIDTH(32)
) inst0 (
    .out(inst0_out)
);
wire _guard0 = 1;
assign p2 = inst0_out;
// COMPONENT END: comp47
endmodule
module comp49(
  output logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp49
logic [31:0] inst0_p2;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_p2;
logic inst1_clk;
logic inst1_reset;
logic [31:0] inst2_p2;
logic inst2_reset;
logic inst2_clk;
logic [31:0] inst3_p4;
logic inst3_clk;
logic inst3_reset;
logic [31:0] inst4_p2;
logic inst4_clk;
logic inst4_reset;
logic [31:0] inst5_p4;
logic inst5_clk;
logic inst5_reset;
logic [31:0] inst6_p2;
logic inst6_reset;
logic inst6_clk;
logic [31:0] inst7_p4;
logic inst7_reset;
logic inst7_clk;
logic [31:0] inst8_p2;
logic inst8_reset;
logic inst8_clk;
logic [31:0] inst9_p4;
logic inst9_reset;
logic inst9_clk;
logic [31:0] inst10_p4;
logic inst10_clk;
logic inst10_reset;
logic [31:0] inst11_p4;
logic inst11_reset;
logic inst11_clk;
logic [31:0] inst12_p4;
logic inst12_clk;
logic inst12_reset;
logic [31:0] inst13_p4;
logic inst13_clk;
logic inst13_reset;
logic [31:0] inst14_p4;
logic inst14_reset;
logic inst14_clk;
logic [31:0] inst15_p4;
logic inst15_clk;
logic inst15_reset;
comp38 inst0 (
    .clk(inst0_clk),
    .p2(inst0_p2),
    .reset(inst0_reset)
);
comp39 inst1 (
    .clk(inst1_clk),
    .p2(inst1_p2),
    .reset(inst1_reset)
);
comp40 inst2 (
    .clk(inst2_clk),
    .p2(inst2_p2),
    .reset(inst2_reset)
);
comp42 inst3 (
    .clk(inst3_clk),
    .p4(inst3_p4),
    .reset(inst3_reset)
);
comp43 inst4 (
    .clk(inst4_clk),
    .p2(inst4_p2),
    .reset(inst4_reset)
);
comp44 inst5 (
    .clk(inst5_clk),
    .p4(inst5_p4),
    .reset(inst5_reset)
);
comp45 inst6 (
    .clk(inst6_clk),
    .p2(inst6_p2),
    .reset(inst6_reset)
);
comp46 inst7 (
    .clk(inst7_clk),
    .p4(inst7_p4),
    .reset(inst7_reset)
);
comp47 inst8 (
    .clk(inst8_clk),
    .p2(inst8_p2),
    .reset(inst8_reset)
);
comp48 inst9 (
    .clk(inst9_clk),
    .p4(inst9_p4),
    .reset(inst9_reset)
);
comp42 inst10 (
    .clk(inst10_clk),
    .p4(inst10_p4),
    .reset(inst10_reset)
);
comp46 inst11 (
    .clk(inst11_clk),
    .p4(inst11_p4),
    .reset(inst11_reset)
);
comp44 inst12 (
    .clk(inst12_clk),
    .p4(inst12_p4),
    .reset(inst12_reset)
);
comp44 inst13 (
    .clk(inst13_clk),
    .p4(inst13_p4),
    .reset(inst13_reset)
);
comp46 inst14 (
    .clk(inst14_clk),
    .p4(inst14_p4),
    .reset(inst14_reset)
);
comp42 inst15 (
    .clk(inst15_clk),
    .p4(inst15_p4),
    .reset(inst15_reset)
);
wire _guard0 = 1;
assign p19 = inst2_p2;
assign p28 = inst11_p4;
assign p29 = inst12_p4;
assign p17 = inst0_p2;
assign p20 = inst3_p4;
assign p21 = inst4_p2;
assign p23 = inst6_p2;
assign p25 = inst8_p2;
assign p18 = inst1_p2;
assign p30 = inst13_p4;
assign p24 = inst7_p4;
assign p32 = inst15_p4;
assign p26 = inst9_p4;
assign p31 = inst14_p4;
assign p27 = inst10_p4;
assign p22 = inst5_p4;
assign inst5_clk = clk;
assign inst5_reset = reset;
assign inst15_clk = clk;
assign inst15_reset = reset;
assign inst8_clk = clk;
assign inst8_reset = reset;
assign inst12_clk = clk;
assign inst12_reset = reset;
assign inst3_clk = clk;
assign inst3_reset = reset;
assign inst9_clk = clk;
assign inst9_reset = reset;
assign inst1_clk = clk;
assign inst1_reset = reset;
assign inst0_clk = clk;
assign inst0_reset = reset;
assign inst7_clk = clk;
assign inst7_reset = reset;
assign inst6_clk = clk;
assign inst6_reset = reset;
assign inst14_clk = clk;
assign inst14_reset = reset;
assign inst2_clk = clk;
assign inst2_reset = reset;
assign inst4_clk = clk;
assign inst4_reset = reset;
assign inst10_clk = clk;
assign inst10_reset = reset;
assign inst11_clk = clk;
assign inst11_reset = reset;
assign inst13_clk = clk;
assign inst13_reset = reset;
// COMPONENT END: comp49
endmodule
module comp53(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp53
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p10;
assign p29 = p11;
assign p20 = p2;
assign p21 = p3;
assign p23 = p3;
assign p25 = p3;
assign p18 = p2;
assign p30 = p10;
assign p24 = p2;
assign p32 = p10;
assign p26 = p10;
assign p31 = p11;
assign p27 = p11;
assign p33 = p11;
assign p22 = p2;
// COMPONENT END: comp53
endmodule
module comp55(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp55
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p12;
assign p29 = p13;
assign p20 = p4;
assign p21 = p5;
assign p23 = p7;
assign p25 = p9;
assign p18 = p2;
assign p30 = p14;
assign p24 = p8;
assign p32 = p16;
assign p26 = p10;
assign p31 = p15;
assign p27 = p11;
assign p33 = p17;
assign p22 = p6;
// COMPONENT END: comp55
endmodule
module comp50(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  output logic [31:0] p40,
  output logic [31:0] p41,
  output logic [31:0] p42,
  output logic [31:0] p43,
  output logic [31:0] p44,
  output logic [31:0] p45,
  output logic [31:0] p46,
  output logic [31:0] p47,
  output logic [31:0] p48,
  output logic [31:0] p49,
  output logic [31:0] p50,
  output logic [31:0] p51,
  output logic [31:0] p52,
  output logic [31:0] p53,
  output logic [31:0] p54,
  output logic [31:0] p55,
  output logic [31:0] p56,
  output logic [31:0] p57,
  output logic [31:0] p58,
  output logic [31:0] p59,
  output logic [31:0] p60,
  output logic [31:0] p61,
  output logic [31:0] p62,
  output logic [31:0] p63,
  output logic [31:0] p64,
  output logic [31:0] p65,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp50
wire _guard0 = 1;
assign p38 = p10;
assign p40 = p26;
assign p47 = p15;
assign p65 = p33;
assign p52 = p20;
assign p59 = p9;
assign p56 = p28;
assign p60 = p24;
assign p64 = p32;
assign p36 = p18;
assign p39 = p11;
assign p46 = p14;
assign p51 = p5;
assign p54 = p12;
assign p45 = p23;
assign p53 = p21;
assign p58 = p8;
assign p50 = p4;
assign p41 = p27;
assign p43 = p7;
assign p63 = p17;
assign p42 = p6;
assign p48 = p30;
assign p49 = p31;
assign p61 = p25;
assign p62 = p16;
assign p34 = p2;
assign p35 = p3;
assign p57 = p29;
assign p37 = p19;
assign p44 = p22;
assign p55 = p13;
// COMPONENT END: comp50
endmodule
module comp54(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp54
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p10;
assign p29 = p11;
assign p20 = p2;
assign p21 = p3;
assign p23 = p7;
assign p25 = p7;
assign p18 = p2;
assign p30 = p14;
assign p24 = p6;
assign p32 = p14;
assign p26 = p10;
assign p31 = p15;
assign p27 = p11;
assign p33 = p15;
assign p22 = p6;
// COMPONENT END: comp54
endmodule
module comp34(
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp34
logic [31:0] inst0_in0_r;
logic [31:0] inst0_in0_i;
logic [31:0] inst0_in1_r;
logic [31:0] inst0_in1_i;
logic [31:0] inst0_twd_r;
logic [31:0] inst0_twd_i;
logic [127:0] inst0_out;
logic inst0_clk;
logic [127:0] inst1_in;
logic [31:0] inst1_out;
logic [127:0] inst2_in;
logic [31:0] inst2_out;
logic [127:0] inst3_in;
logic [31:0] inst3_out;
logic [127:0] inst4_in;
logic [31:0] inst4_out;
Butterfly_Exp8_Mant23 inst0 (
    .clk(inst0_clk),
    .in0_i(inst0_in0_i),
    .in0_r(inst0_in0_r),
    .in1_i(inst0_in1_i),
    .in1_r(inst0_in1_r),
    .out(inst0_out),
    .twd_i(inst0_twd_i),
    .twd_r(inst0_twd_r)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(96),
    .MSB(127),
    .OUT_WIDTH(32)
) inst1 (
    .in(inst1_in),
    .out(inst1_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(64),
    .MSB(95),
    .OUT_WIDTH(32)
) inst2 (
    .in(inst2_in),
    .out(inst2_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(32),
    .MSB(63),
    .OUT_WIDTH(32)
) inst3 (
    .in(inst3_in),
    .out(inst3_out)
);
Slice # (
    .IN_WIDTH(128),
    .LSB(0),
    .MSB(31),
    .OUT_WIDTH(32)
) inst4 (
    .in(inst4_in),
    .out(inst4_out)
);
wire _guard0 = 1;
assign p28 = inst3_out;
assign p29 = inst4_out;
assign p26 = inst1_out;
assign p27 = inst2_out;
assign inst3_in = inst0_out;
assign inst1_in = inst0_out;
assign inst0_in1_i = p23;
assign inst0_twd_i = p25;
assign inst0_clk = clk;
assign inst0_in0_i = p21;
assign inst0_in1_r = p22;
assign inst0_twd_r = p24;
assign inst0_in0_r = p20;
assign inst2_in = inst0_out;
assign inst4_in = inst0_out;
// COMPONENT END: comp34
endmodule
module comp91(
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  output logic [1023:0] p37,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp91
logic [31:0] inst0_p7;
logic [31:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [31:0] inst0_p38;
logic [1023:0] inst0_p39;
logic inst0_reset;
logic inst0_clk;
comp90 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p39(inst0_p39),
    .p7(inst0_p7),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
wire _guard0 = 1;
assign p37 = inst0_p39;
assign inst0_p19 = p17;
assign inst0_p28 = p26;
assign inst0_p29 = p27;
assign inst0_p38 = p36;
assign inst0_p12 = p10;
assign inst0_p16 = p14;
assign inst0_p9 = p7;
assign inst0_p15 = p13;
assign inst0_p17 = p15;
assign inst0_p20 = p18;
assign inst0_p21 = p19;
assign inst0_p23 = p21;
assign inst0_clk = clk;
assign inst0_p11 = p9;
assign inst0_p25 = p23;
assign inst0_p36 = p34;
assign inst0_p8 = p6;
assign inst0_p10 = p8;
assign inst0_reset = reset;
assign inst0_p13 = p11;
assign inst0_p18 = p16;
assign inst0_p30 = p28;
assign inst0_p7 = p5;
assign inst0_p24 = p22;
assign inst0_p32 = p30;
assign inst0_p14 = p12;
assign inst0_p26 = p24;
assign inst0_p31 = p29;
assign inst0_p27 = p25;
assign inst0_p33 = p31;
assign inst0_p22 = p20;
assign inst0_p34 = p32;
assign inst0_p35 = p33;
assign inst0_p37 = p35;
// COMPONENT END: comp91
endmodule
module comp36(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  output logic [31:0] p34,
  output logic [31:0] p35,
  output logic [31:0] p36,
  output logic [31:0] p37,
  output logic [31:0] p38,
  output logic [31:0] p39,
  output logic [31:0] p40,
  output logic [31:0] p41,
  output logic [31:0] p42,
  output logic [31:0] p43,
  output logic [31:0] p44,
  output logic [31:0] p45,
  output logic [31:0] p46,
  output logic [31:0] p47,
  output logic [31:0] p48,
  output logic [31:0] p49,
  output logic [31:0] p50,
  output logic [31:0] p51,
  output logic [31:0] p52,
  output logic [31:0] p53,
  output logic [31:0] p54,
  output logic [31:0] p55,
  output logic [31:0] p56,
  output logic [31:0] p57,
  output logic [31:0] p58,
  output logic [31:0] p59,
  output logic [31:0] p60,
  output logic [31:0] p61,
  output logic [31:0] p62,
  output logic [31:0] p63,
  output logic [31:0] p64,
  output logic [31:0] p65,
  input logic reset,
  input logic clk
);
// COMPONENT START: comp36
wire _guard0 = 1;
assign p38 = p10;
assign p40 = p14;
assign p47 = p27;
assign p65 = p33;
assign p52 = p8;
assign p59 = p21;
assign p56 = p16;
assign p60 = p24;
assign p64 = p32;
assign p36 = p6;
assign p39 = p11;
assign p46 = p26;
assign p51 = p5;
assign p54 = p12;
assign p45 = p23;
assign p53 = p9;
assign p58 = p20;
assign p50 = p4;
assign p41 = p15;
assign p43 = p19;
assign p63 = p29;
assign p42 = p18;
assign p48 = p30;
assign p49 = p31;
assign p61 = p25;
assign p62 = p28;
assign p34 = p2;
assign p35 = p3;
assign p57 = p17;
assign p37 = p7;
assign p44 = p22;
assign p55 = p13;
// COMPONENT END: comp36
endmodule
module comp52(
  input logic [31:0] p2,
  input logic [31:0] p3,
  input logic [31:0] p4,
  input logic [31:0] p5,
  input logic [31:0] p6,
  input logic [31:0] p7,
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  output logic [31:0] p18,
  output logic [31:0] p19,
  output logic [31:0] p20,
  output logic [31:0] p21,
  output logic [31:0] p22,
  output logic [31:0] p23,
  output logic [31:0] p24,
  output logic [31:0] p25,
  output logic [31:0] p26,
  output logic [31:0] p27,
  output logic [31:0] p28,
  output logic [31:0] p29,
  output logic [31:0] p30,
  output logic [31:0] p31,
  output logic [31:0] p32,
  output logic [31:0] p33,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp52
wire _guard0 = 1;
assign p19 = p3;
assign p28 = p2;
assign p29 = p3;
assign p20 = p2;
assign p21 = p3;
assign p23 = p3;
assign p25 = p3;
assign p18 = p2;
assign p30 = p2;
assign p24 = p2;
assign p32 = p2;
assign p26 = p2;
assign p31 = p3;
assign p27 = p3;
assign p33 = p3;
assign p22 = p2;
// COMPONENT END: comp52
endmodule
module comp35(
  input logic [31:0] p43,
  input logic [31:0] p44,
  input logic [31:0] p45,
  input logic [31:0] p46,
  input logic [31:0] p47,
  input logic [31:0] p48,
  input logic [31:0] p49,
  input logic [31:0] p50,
  input logic [31:0] p51,
  input logic [31:0] p52,
  input logic [31:0] p53,
  input logic [31:0] p54,
  input logic [31:0] p55,
  input logic [31:0] p56,
  input logic [31:0] p57,
  input logic [31:0] p58,
  input logic [31:0] p59,
  input logic [31:0] p60,
  input logic [31:0] p61,
  input logic [31:0] p62,
  input logic [31:0] p63,
  input logic [31:0] p64,
  input logic [31:0] p65,
  input logic [31:0] p66,
  input logic [31:0] p67,
  input logic [31:0] p68,
  input logic [31:0] p69,
  input logic [31:0] p70,
  input logic [31:0] p71,
  input logic [31:0] p72,
  input logic [31:0] p73,
  input logic [31:0] p74,
  input logic [31:0] p75,
  input logic [31:0] p76,
  input logic [31:0] p77,
  input logic [31:0] p78,
  input logic [31:0] p79,
  input logic [31:0] p80,
  input logic [31:0] p81,
  input logic [31:0] p82,
  input logic [31:0] p83,
  input logic [31:0] p84,
  input logic [31:0] p85,
  input logic [31:0] p86,
  input logic [31:0] p87,
  input logic [31:0] p88,
  input logic [31:0] p89,
  input logic [31:0] p90,
  output logic [31:0] p91,
  output logic [31:0] p92,
  output logic [31:0] p93,
  output logic [31:0] p94,
  output logic [31:0] p95,
  output logic [31:0] p96,
  output logic [31:0] p97,
  output logic [31:0] p98,
  output logic [31:0] p99,
  output logic [31:0] p100,
  output logic [31:0] p101,
  output logic [31:0] p102,
  output logic [31:0] p103,
  output logic [31:0] p104,
  output logic [31:0] p105,
  output logic [31:0] p106,
  output logic [31:0] p107,
  output logic [31:0] p108,
  output logic [31:0] p109,
  output logic [31:0] p110,
  output logic [31:0] p111,
  output logic [31:0] p112,
  output logic [31:0] p113,
  output logic [31:0] p114,
  output logic [31:0] p115,
  output logic [31:0] p116,
  output logic [31:0] p117,
  output logic [31:0] p118,
  output logic [31:0] p119,
  output logic [31:0] p120,
  output logic [31:0] p121,
  output logic [31:0] p122,
  input logic ev0,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp35
logic ev00__0;
logic ev00__1;
logic ev00__2;
logic ev00__3;
logic ev00__4;
logic ev00__5;
logic ev00__6;
logic ev00__7;
logic ev00__8;
logic ev00__9;
logic ev00__10;
logic ev00__11;
logic ev00__12;
logic ev00__13;
logic ev00__14;
logic ev00__15;
logic ev00__16;
logic ev00__17;
logic ev00__18;
logic ev00__19;
logic ev00__20;
logic ev00__21;
logic ev00__22;
logic ev00__23;
logic ev00__24;
logic ev00__25;
logic ev00__26;
logic ev00__27;
logic ev00__28;
logic ev00__29;
logic ev00__30;
logic ev00_clk;
logic ev00_reset;
logic ev00_go;
logic ev00_done;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic inst1_clk;
logic inst1_reset;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic inst2_clk;
logic inst2_reset;
logic [31:0] inst3_p20;
logic [31:0] inst3_p21;
logic [31:0] inst3_p22;
logic [31:0] inst3_p23;
logic [31:0] inst3_p24;
logic [31:0] inst3_p25;
logic [31:0] inst3_p26;
logic [31:0] inst3_p27;
logic [31:0] inst3_p28;
logic [31:0] inst3_p29;
logic inst3_clk;
logic inst3_reset;
logic [31:0] inst4_p20;
logic [31:0] inst4_p21;
logic [31:0] inst4_p22;
logic [31:0] inst4_p23;
logic [31:0] inst4_p24;
logic [31:0] inst4_p25;
logic [31:0] inst4_p26;
logic [31:0] inst4_p27;
logic [31:0] inst4_p28;
logic [31:0] inst4_p29;
logic inst4_clk;
logic inst4_reset;
logic [31:0] inst5_p20;
logic [31:0] inst5_p21;
logic [31:0] inst5_p22;
logic [31:0] inst5_p23;
logic [31:0] inst5_p24;
logic [31:0] inst5_p25;
logic [31:0] inst5_p26;
logic [31:0] inst5_p27;
logic [31:0] inst5_p28;
logic [31:0] inst5_p29;
logic inst5_clk;
logic inst5_reset;
logic [31:0] inst6_p20;
logic [31:0] inst6_p21;
logic [31:0] inst6_p22;
logic [31:0] inst6_p23;
logic [31:0] inst6_p24;
logic [31:0] inst6_p25;
logic [31:0] inst6_p26;
logic [31:0] inst6_p27;
logic [31:0] inst6_p28;
logic [31:0] inst6_p29;
logic inst6_clk;
logic inst6_reset;
logic [31:0] inst7_p20;
logic [31:0] inst7_p21;
logic [31:0] inst7_p22;
logic [31:0] inst7_p23;
logic [31:0] inst7_p24;
logic [31:0] inst7_p25;
logic [31:0] inst7_p26;
logic [31:0] inst7_p27;
logic [31:0] inst7_p28;
logic [31:0] inst7_p29;
logic inst7_clk;
logic inst7_reset;
logic [31:0] inst8_p20;
logic [31:0] inst8_p21;
logic [31:0] inst8_p22;
logic [31:0] inst8_p23;
logic [31:0] inst8_p24;
logic [31:0] inst8_p25;
logic [31:0] inst8_p26;
logic [31:0] inst8_p27;
logic [31:0] inst8_p28;
logic [31:0] inst8_p29;
logic inst8_clk;
logic inst8_reset;
fsm_31 ev00 (
    ._0(ev00__0),
    ._1(ev00__1),
    ._10(ev00__10),
    ._11(ev00__11),
    ._12(ev00__12),
    ._13(ev00__13),
    ._14(ev00__14),
    ._15(ev00__15),
    ._16(ev00__16),
    ._17(ev00__17),
    ._18(ev00__18),
    ._19(ev00__19),
    ._2(ev00__2),
    ._20(ev00__20),
    ._21(ev00__21),
    ._22(ev00__22),
    ._23(ev00__23),
    ._24(ev00__24),
    ._25(ev00__25),
    ._26(ev00__26),
    ._27(ev00__27),
    ._28(ev00__28),
    ._29(ev00__29),
    ._3(ev00__3),
    ._30(ev00__30),
    ._4(ev00__4),
    ._5(ev00__5),
    ._6(ev00__6),
    ._7(ev00__7),
    ._8(ev00__8),
    ._9(ev00__9),
    .clk(ev00_clk),
    .done(ev00_done),
    .go(ev00_go),
    .reset(ev00_reset)
);
comp34 inst1 (
    .clk(inst1_clk),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .reset(inst1_reset)
);
comp34 inst2 (
    .clk(inst2_clk),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .reset(inst2_reset)
);
comp34 inst3 (
    .clk(inst3_clk),
    .p20(inst3_p20),
    .p21(inst3_p21),
    .p22(inst3_p22),
    .p23(inst3_p23),
    .p24(inst3_p24),
    .p25(inst3_p25),
    .p26(inst3_p26),
    .p27(inst3_p27),
    .p28(inst3_p28),
    .p29(inst3_p29),
    .reset(inst3_reset)
);
comp34 inst4 (
    .clk(inst4_clk),
    .p20(inst4_p20),
    .p21(inst4_p21),
    .p22(inst4_p22),
    .p23(inst4_p23),
    .p24(inst4_p24),
    .p25(inst4_p25),
    .p26(inst4_p26),
    .p27(inst4_p27),
    .p28(inst4_p28),
    .p29(inst4_p29),
    .reset(inst4_reset)
);
comp34 inst5 (
    .clk(inst5_clk),
    .p20(inst5_p20),
    .p21(inst5_p21),
    .p22(inst5_p22),
    .p23(inst5_p23),
    .p24(inst5_p24),
    .p25(inst5_p25),
    .p26(inst5_p26),
    .p27(inst5_p27),
    .p28(inst5_p28),
    .p29(inst5_p29),
    .reset(inst5_reset)
);
comp34 inst6 (
    .clk(inst6_clk),
    .p20(inst6_p20),
    .p21(inst6_p21),
    .p22(inst6_p22),
    .p23(inst6_p23),
    .p24(inst6_p24),
    .p25(inst6_p25),
    .p26(inst6_p26),
    .p27(inst6_p27),
    .p28(inst6_p28),
    .p29(inst6_p29),
    .reset(inst6_reset)
);
comp34 inst7 (
    .clk(inst7_clk),
    .p20(inst7_p20),
    .p21(inst7_p21),
    .p22(inst7_p22),
    .p23(inst7_p23),
    .p24(inst7_p24),
    .p25(inst7_p25),
    .p26(inst7_p26),
    .p27(inst7_p27),
    .p28(inst7_p28),
    .p29(inst7_p29),
    .reset(inst7_reset)
);
comp34 inst8 (
    .clk(inst8_clk),
    .p20(inst8_p20),
    .p21(inst8_p21),
    .p22(inst8_p22),
    .p23(inst8_p23),
    .p24(inst8_p24),
    .p25(inst8_p25),
    .p26(inst8_p26),
    .p27(inst8_p27),
    .p28(inst8_p28),
    .p29(inst8_p29),
    .reset(inst8_reset)
);
wire _guard0 = 1;
wire _guard1 = ev00__30;
wire _guard2 = ev00__30;
wire _guard3 = ev00__30;
wire _guard4 = ev00__30;
wire _guard5 = ev00__30;
wire _guard6 = ev00__30;
wire _guard7 = ev00__30;
wire _guard8 = ev00__30;
wire _guard9 = ev00__30;
wire _guard10 = ev00__30;
wire _guard11 = ev00__30;
wire _guard12 = ev00__30;
wire _guard13 = ev00__30;
wire _guard14 = ev00__30;
wire _guard15 = ev00__30;
wire _guard16 = ev00__30;
wire _guard17 = ev00__30;
wire _guard18 = ev00__30;
wire _guard19 = ev00__30;
wire _guard20 = ev00__30;
wire _guard21 = ev00__30;
wire _guard22 = ev00__30;
wire _guard23 = ev00__30;
wire _guard24 = ev00__30;
wire _guard25 = ev00__30;
wire _guard26 = ev00__30;
wire _guard27 = ev00__30;
wire _guard28 = ev00__30;
wire _guard29 = ev00__30;
wire _guard30 = ev00__30;
wire _guard31 = ev00__30;
wire _guard32 = ev00__30;
wire _guard33 = ev00__0;
wire _guard34 = ev00__0;
wire _guard35 = ev00__0;
wire _guard36 = ev00__0;
wire _guard37 = ev00__0;
wire _guard38 = ev00__0;
wire _guard39 = ev00__0;
wire _guard40 = ev00__0;
wire _guard41 = ev00__0;
wire _guard42 = ev00__0;
wire _guard43 = ev00__0;
wire _guard44 = ev00__0;
wire _guard45 = ev00__0;
wire _guard46 = ev00__0;
wire _guard47 = ev00__0;
wire _guard48 = ev00__0;
wire _guard49 = ev00__0;
wire _guard50 = ev00__0;
wire _guard51 = ev00__0;
wire _guard52 = ev00__0;
wire _guard53 = ev00__0;
wire _guard54 = ev00__0;
wire _guard55 = ev00__0;
wire _guard56 = ev00__0;
wire _guard57 = ev00__0;
wire _guard58 = ev00__0;
wire _guard59 = ev00__0;
wire _guard60 = ev00__0;
wire _guard61 = ev00__0;
wire _guard62 = ev00__0;
wire _guard63 = ev00__0;
wire _guard64 = ev00__0;
wire _guard65 = ev00__0;
wire _guard66 = ev00__0;
wire _guard67 = ev00__0;
wire _guard68 = ev00__0;
wire _guard69 = ev00__0;
wire _guard70 = ev00__0;
wire _guard71 = ev00__0;
wire _guard72 = ev00__0;
wire _guard73 = ev00__0;
wire _guard74 = ev00__0;
wire _guard75 = ev00__0;
wire _guard76 = ev00__0;
wire _guard77 = ev00__0;
wire _guard78 = ev00__0;
wire _guard79 = ev00__0;
wire _guard80 = ev00__0;
assign p104 =
  _guard1 ? inst4_p27 :
  32'd0;
assign p120 =
  _guard2 ? inst8_p27 :
  32'd0;
assign p110 =
  _guard3 ? inst5_p29 :
  32'd0;
assign p115 =
  _guard4 ? inst7_p26 :
  32'd0;
assign p116 =
  _guard5 ? inst7_p27 :
  32'd0;
assign p121 =
  _guard6 ? inst8_p28 :
  32'd0;
assign p94 =
  _guard7 ? inst1_p29 :
  32'd0;
assign p99 =
  _guard8 ? inst3_p26 :
  32'd0;
assign p102 =
  _guard9 ? inst3_p29 :
  32'd0;
assign p98 =
  _guard10 ? inst2_p29 :
  32'd0;
assign p107 =
  _guard11 ? inst5_p26 :
  32'd0;
assign p109 =
  _guard12 ? inst5_p28 :
  32'd0;
assign p111 =
  _guard13 ? inst6_p26 :
  32'd0;
assign p96 =
  _guard14 ? inst2_p27 :
  32'd0;
assign p100 =
  _guard15 ? inst3_p27 :
  32'd0;
assign p113 =
  _guard16 ? inst6_p28 :
  32'd0;
assign p117 =
  _guard17 ? inst7_p28 :
  32'd0;
assign p119 =
  _guard18 ? inst8_p26 :
  32'd0;
assign p97 =
  _guard19 ? inst2_p28 :
  32'd0;
assign p112 =
  _guard20 ? inst6_p27 :
  32'd0;
assign p92 =
  _guard21 ? inst1_p27 :
  32'd0;
assign p108 =
  _guard22 ? inst5_p27 :
  32'd0;
assign p103 =
  _guard23 ? inst4_p26 :
  32'd0;
assign p105 =
  _guard24 ? inst4_p28 :
  32'd0;
assign p114 =
  _guard25 ? inst6_p29 :
  32'd0;
assign p118 =
  _guard26 ? inst7_p29 :
  32'd0;
assign p93 =
  _guard27 ? inst1_p28 :
  32'd0;
assign p95 =
  _guard28 ? inst2_p26 :
  32'd0;
assign p106 =
  _guard29 ? inst4_p29 :
  32'd0;
assign p91 =
  _guard30 ? inst1_p26 :
  32'd0;
assign p101 =
  _guard31 ? inst3_p28 :
  32'd0;
assign p122 =
  _guard32 ? inst8_p29 :
  32'd0;
assign inst5_p20 = p59;
assign inst5_p21 = p60;
assign inst5_p23 = p62;
assign inst5_clk = clk;
assign inst5_p25 = p84;
assign inst5_reset = reset;
assign inst5_p24 = p83;
assign inst5_p22 = p61;
assign inst8_p20 = p71;
assign inst8_p21 = p72;
assign inst8_p23 = p74;
assign inst8_clk = clk;
assign inst8_p25 = p90;
assign inst8_reset = reset;
assign inst8_p24 = p89;
assign inst8_p22 = p73;
assign inst3_p20 = p51;
assign inst3_p21 = p52;
assign inst3_p23 = p54;
assign inst3_clk = clk;
assign inst3_p25 = p80;
assign inst3_reset = reset;
assign inst3_p24 = p79;
assign inst3_p22 = p53;
assign inst1_p20 = p43;
assign inst1_p21 = p44;
assign inst1_p23 = p46;
assign inst1_clk = clk;
assign inst1_p25 = p76;
assign inst1_reset = reset;
assign inst1_p24 = p75;
assign inst1_p22 = p45;
assign inst7_p20 = p67;
assign inst7_p21 = p68;
assign inst7_p23 = p70;
assign inst7_clk = clk;
assign inst7_p25 = p88;
assign inst7_reset = reset;
assign inst7_p24 = p87;
assign inst7_p22 = p69;
assign ev00_clk = clk;
assign ev00_go = ev0;
assign ev00_reset = reset;
assign inst6_p20 = p63;
assign inst6_p21 = p64;
assign inst6_p23 = p66;
assign inst6_clk = clk;
assign inst6_p25 = p86;
assign inst6_reset = reset;
assign inst6_p24 = p85;
assign inst6_p22 = p65;
assign inst2_p20 = p47;
assign inst2_p21 = p48;
assign inst2_p23 = p50;
assign inst2_clk = clk;
assign inst2_p25 = p78;
assign inst2_reset = reset;
assign inst2_p24 = p77;
assign inst2_p22 = p49;
assign inst4_p20 = p55;
assign inst4_p21 = p56;
assign inst4_p23 = p58;
assign inst4_clk = clk;
assign inst4_p25 = p82;
assign inst4_reset = reset;
assign inst4_p24 = p81;
assign inst4_p22 = p57;
// COMPONENT END: comp35
endmodule
module comp92(
  input logic [31:0] p108,
  input logic [31:0] p109,
  input logic [31:0] p110,
  input logic [31:0] p111,
  input logic [31:0] p112,
  input logic [31:0] p113,
  input logic [31:0] p114,
  input logic [31:0] p115,
  input logic [31:0] p116,
  input logic [31:0] p117,
  input logic [31:0] p118,
  input logic [31:0] p119,
  input logic [31:0] p120,
  input logic [31:0] p121,
  input logic [31:0] p122,
  input logic [31:0] p123,
  input logic [31:0] p124,
  input logic [31:0] p125,
  input logic [31:0] p126,
  input logic [31:0] p127,
  input logic [31:0] p128,
  input logic [31:0] p129,
  input logic [31:0] p130,
  input logic [31:0] p131,
  input logic [31:0] p132,
  input logic [31:0] p133,
  input logic [31:0] p134,
  input logic [31:0] p135,
  input logic [31:0] p136,
  input logic [31:0] p137,
  input logic [31:0] p138,
  input logic [31:0] p139,
  output logic [31:0] p140,
  output logic [31:0] p141,
  output logic [31:0] p142,
  output logic [31:0] p143,
  output logic [31:0] p144,
  output logic [31:0] p145,
  output logic [31:0] p146,
  output logic [31:0] p147,
  output logic [31:0] p148,
  output logic [31:0] p149,
  output logic [31:0] p150,
  output logic [31:0] p151,
  output logic [31:0] p152,
  output logic [31:0] p153,
  output logic [31:0] p154,
  output logic [31:0] p155,
  output logic [31:0] p156,
  output logic [31:0] p157,
  output logic [31:0] p158,
  output logic [31:0] p159,
  output logic [31:0] p160,
  output logic [31:0] p161,
  output logic [31:0] p162,
  output logic [31:0] p163,
  output logic [31:0] p164,
  output logic [31:0] p165,
  output logic [31:0] p166,
  output logic [31:0] p167,
  output logic [31:0] p168,
  output logic [31:0] p169,
  output logic [31:0] p170,
  output logic [31:0] p171,
  input logic ev0,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp92
logic [6:0] ev00__0state;
logic ev00__0_0;
logic [6:0] ev00__1state;
logic ev00__1_0;
logic ev00_clk;
logic ev00_reset;
logic ev00_go;
logic ev00_done;
logic [31:0] inst0_p43;
logic [31:0] inst0_p44;
logic [31:0] inst0_p45;
logic [31:0] inst0_p46;
logic [31:0] inst0_p47;
logic [31:0] inst0_p48;
logic [31:0] inst0_p49;
logic [31:0] inst0_p50;
logic [31:0] inst0_p51;
logic [31:0] inst0_p52;
logic [31:0] inst0_p53;
logic [31:0] inst0_p54;
logic [31:0] inst0_p55;
logic [31:0] inst0_p56;
logic [31:0] inst0_p57;
logic [31:0] inst0_p58;
logic [31:0] inst0_p59;
logic [31:0] inst0_p60;
logic [31:0] inst0_p61;
logic [31:0] inst0_p62;
logic [31:0] inst0_p63;
logic [31:0] inst0_p64;
logic [31:0] inst0_p65;
logic [31:0] inst0_p66;
logic [31:0] inst0_p67;
logic [31:0] inst0_p68;
logic [31:0] inst0_p69;
logic [31:0] inst0_p70;
logic [31:0] inst0_p71;
logic [31:0] inst0_p72;
logic [31:0] inst0_p73;
logic [31:0] inst0_p74;
logic [31:0] inst0_p75;
logic [31:0] inst0_p76;
logic [31:0] inst0_p77;
logic [31:0] inst0_p78;
logic [31:0] inst0_p79;
logic [31:0] inst0_p80;
logic [31:0] inst0_p81;
logic [31:0] inst0_p82;
logic [31:0] inst0_p83;
logic [31:0] inst0_p84;
logic [31:0] inst0_p85;
logic [31:0] inst0_p86;
logic [31:0] inst0_p87;
logic [31:0] inst0_p88;
logic [31:0] inst0_p89;
logic [31:0] inst0_p90;
logic [31:0] inst0_p91;
logic [31:0] inst0_p92;
logic [31:0] inst0_p93;
logic [31:0] inst0_p94;
logic [31:0] inst0_p95;
logic [31:0] inst0_p96;
logic [31:0] inst0_p97;
logic [31:0] inst0_p98;
logic [31:0] inst0_p99;
logic [31:0] inst0_p100;
logic [31:0] inst0_p101;
logic [31:0] inst0_p102;
logic [31:0] inst0_p103;
logic [31:0] inst0_p104;
logic [31:0] inst0_p105;
logic [31:0] inst0_p106;
logic [31:0] inst0_p107;
logic [31:0] inst0_p108;
logic [31:0] inst0_p109;
logic [31:0] inst0_p110;
logic [31:0] inst0_p111;
logic [31:0] inst0_p112;
logic [31:0] inst0_p113;
logic [31:0] inst0_p114;
logic [31:0] inst0_p115;
logic [31:0] inst0_p116;
logic [31:0] inst0_p117;
logic [31:0] inst0_p118;
logic [31:0] inst0_p119;
logic [31:0] inst0_p120;
logic [31:0] inst0_p121;
logic [31:0] inst0_p122;
logic inst0_ev0;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_p2;
logic [31:0] inst1_p3;
logic [31:0] inst1_p4;
logic [31:0] inst1_p5;
logic [31:0] inst1_p6;
logic [31:0] inst1_p7;
logic [31:0] inst1_p8;
logic [31:0] inst1_p9;
logic [31:0] inst1_p10;
logic [31:0] inst1_p11;
logic [31:0] inst1_p12;
logic [31:0] inst1_p13;
logic [31:0] inst1_p14;
logic [31:0] inst1_p15;
logic [31:0] inst1_p16;
logic [31:0] inst1_p17;
logic [31:0] inst1_p18;
logic [31:0] inst1_p19;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic [31:0] inst1_p30;
logic [31:0] inst1_p31;
logic [31:0] inst1_p32;
logic [31:0] inst1_p33;
logic [31:0] inst1_p34;
logic [31:0] inst1_p35;
logic [31:0] inst1_p36;
logic [31:0] inst1_p37;
logic [31:0] inst1_p38;
logic [31:0] inst1_p39;
logic [31:0] inst1_p40;
logic [31:0] inst1_p41;
logic [31:0] inst1_p42;
logic [31:0] inst1_p43;
logic [31:0] inst1_p44;
logic [31:0] inst1_p45;
logic [31:0] inst1_p46;
logic [31:0] inst1_p47;
logic [31:0] inst1_p48;
logic [31:0] inst1_p49;
logic [31:0] inst1_p50;
logic [31:0] inst1_p51;
logic [31:0] inst1_p52;
logic [31:0] inst1_p53;
logic [31:0] inst1_p54;
logic [31:0] inst1_p55;
logic [31:0] inst1_p56;
logic [31:0] inst1_p57;
logic [31:0] inst1_p58;
logic [31:0] inst1_p59;
logic [31:0] inst1_p60;
logic [31:0] inst1_p61;
logic [31:0] inst1_p62;
logic [31:0] inst1_p63;
logic [31:0] inst1_p64;
logic [31:0] inst1_p65;
logic inst1_reset;
logic inst1_clk;
logic [31:0] inst2_p17;
logic [31:0] inst2_p18;
logic [31:0] inst2_p19;
logic [31:0] inst2_p20;
logic [31:0] inst2_p21;
logic [31:0] inst2_p22;
logic [31:0] inst2_p23;
logic [31:0] inst2_p24;
logic [31:0] inst2_p25;
logic [31:0] inst2_p26;
logic [31:0] inst2_p27;
logic [31:0] inst2_p28;
logic [31:0] inst2_p29;
logic [31:0] inst2_p30;
logic [31:0] inst2_p31;
logic [31:0] inst2_p32;
logic inst2_clk;
logic inst2_reset;
logic [31:0] inst3_p2;
logic [31:0] inst3_p3;
logic [31:0] inst3_p4;
logic [31:0] inst3_p5;
logic [31:0] inst3_p6;
logic [31:0] inst3_p7;
logic [31:0] inst3_p8;
logic [31:0] inst3_p9;
logic [31:0] inst3_p10;
logic [31:0] inst3_p11;
logic [31:0] inst3_p12;
logic [31:0] inst3_p13;
logic [31:0] inst3_p14;
logic [31:0] inst3_p15;
logic [31:0] inst3_p16;
logic [31:0] inst3_p17;
logic [31:0] inst3_p18;
logic [31:0] inst3_p19;
logic [31:0] inst3_p20;
logic [31:0] inst3_p21;
logic [31:0] inst3_p22;
logic [31:0] inst3_p23;
logic [31:0] inst3_p24;
logic [31:0] inst3_p25;
logic [31:0] inst3_p26;
logic [31:0] inst3_p27;
logic [31:0] inst3_p28;
logic [31:0] inst3_p29;
logic [31:0] inst3_p30;
logic [31:0] inst3_p31;
logic [31:0] inst3_p32;
logic [31:0] inst3_p33;
logic [31:0] inst3_p34;
logic [31:0] inst3_p35;
logic [31:0] inst3_p36;
logic [31:0] inst3_p37;
logic [31:0] inst3_p38;
logic [31:0] inst3_p39;
logic [31:0] inst3_p40;
logic [31:0] inst3_p41;
logic [31:0] inst3_p42;
logic [31:0] inst3_p43;
logic [31:0] inst3_p44;
logic [31:0] inst3_p45;
logic [31:0] inst3_p46;
logic [31:0] inst3_p47;
logic [31:0] inst3_p48;
logic [31:0] inst3_p49;
logic [31:0] inst3_p50;
logic [31:0] inst3_p51;
logic [31:0] inst3_p52;
logic [31:0] inst3_p53;
logic [31:0] inst3_p54;
logic [31:0] inst3_p55;
logic [31:0] inst3_p56;
logic [31:0] inst3_p57;
logic [31:0] inst3_p58;
logic [31:0] inst3_p59;
logic [31:0] inst3_p60;
logic [31:0] inst3_p61;
logic [31:0] inst3_p62;
logic [31:0] inst3_p63;
logic [31:0] inst3_p64;
logic [31:0] inst3_p65;
logic inst3_clk;
logic inst3_reset;
logic [1023:0] inst4_in;
logic [1023:0] inst4_out;
logic inst4_clk;
logic inst4_reset;
logic [31:0] inst5_p2;
logic [31:0] inst5_p3;
logic [31:0] inst5_p4;
logic [31:0] inst5_p5;
logic [31:0] inst5_p6;
logic [31:0] inst5_p7;
logic [31:0] inst5_p8;
logic [31:0] inst5_p9;
logic [31:0] inst5_p10;
logic [31:0] inst5_p11;
logic [31:0] inst5_p12;
logic [31:0] inst5_p13;
logic [31:0] inst5_p14;
logic [31:0] inst5_p15;
logic [31:0] inst5_p16;
logic [31:0] inst5_p17;
logic [31:0] inst5_p18;
logic [31:0] inst5_p19;
logic [31:0] inst5_p20;
logic [31:0] inst5_p21;
logic [31:0] inst5_p22;
logic [31:0] inst5_p23;
logic [31:0] inst5_p24;
logic [31:0] inst5_p25;
logic [31:0] inst5_p26;
logic [31:0] inst5_p27;
logic [31:0] inst5_p28;
logic [31:0] inst5_p29;
logic [31:0] inst5_p30;
logic [31:0] inst5_p31;
logic [31:0] inst5_p32;
logic [31:0] inst5_p33;
logic inst5_clk;
logic inst5_reset;
logic [31:0] inst6_p2;
logic [31:0] inst6_p3;
logic [31:0] inst6_p4;
logic [31:0] inst6_p5;
logic [31:0] inst6_p6;
logic [31:0] inst6_p7;
logic [31:0] inst6_p8;
logic [31:0] inst6_p9;
logic [31:0] inst6_p10;
logic [31:0] inst6_p11;
logic [31:0] inst6_p12;
logic [31:0] inst6_p13;
logic [31:0] inst6_p14;
logic [31:0] inst6_p15;
logic [31:0] inst6_p16;
logic [31:0] inst6_p17;
logic [31:0] inst6_p18;
logic [31:0] inst6_p19;
logic [31:0] inst6_p20;
logic [31:0] inst6_p21;
logic [31:0] inst6_p22;
logic [31:0] inst6_p23;
logic [31:0] inst6_p24;
logic [31:0] inst6_p25;
logic [31:0] inst6_p26;
logic [31:0] inst6_p27;
logic [31:0] inst6_p28;
logic [31:0] inst6_p29;
logic [31:0] inst6_p30;
logic [31:0] inst6_p31;
logic [31:0] inst6_p32;
logic [31:0] inst6_p33;
logic inst6_clk;
logic inst6_reset;
logic [31:0] inst7_p2;
logic [31:0] inst7_p3;
logic [31:0] inst7_p4;
logic [31:0] inst7_p5;
logic [31:0] inst7_p6;
logic [31:0] inst7_p7;
logic [31:0] inst7_p8;
logic [31:0] inst7_p9;
logic [31:0] inst7_p10;
logic [31:0] inst7_p11;
logic [31:0] inst7_p12;
logic [31:0] inst7_p13;
logic [31:0] inst7_p14;
logic [31:0] inst7_p15;
logic [31:0] inst7_p16;
logic [31:0] inst7_p17;
logic [31:0] inst7_p18;
logic [31:0] inst7_p19;
logic [31:0] inst7_p20;
logic [31:0] inst7_p21;
logic [31:0] inst7_p22;
logic [31:0] inst7_p23;
logic [31:0] inst7_p24;
logic [31:0] inst7_p25;
logic [31:0] inst7_p26;
logic [31:0] inst7_p27;
logic [31:0] inst7_p28;
logic [31:0] inst7_p29;
logic [31:0] inst7_p30;
logic [31:0] inst7_p31;
logic [31:0] inst7_p32;
logic [31:0] inst7_p33;
logic inst7_reset;
logic inst7_clk;
logic [31:0] inst8_p2;
logic [31:0] inst8_p3;
logic [31:0] inst8_p4;
logic [31:0] inst8_p5;
logic [31:0] inst8_p6;
logic [31:0] inst8_p7;
logic [31:0] inst8_p8;
logic [31:0] inst8_p9;
logic [31:0] inst8_p10;
logic [31:0] inst8_p11;
logic [31:0] inst8_p12;
logic [31:0] inst8_p13;
logic [31:0] inst8_p14;
logic [31:0] inst8_p15;
logic [31:0] inst8_p16;
logic [31:0] inst8_p17;
logic [31:0] inst8_p18;
logic [31:0] inst8_p19;
logic [31:0] inst8_p20;
logic [31:0] inst8_p21;
logic [31:0] inst8_p22;
logic [31:0] inst8_p23;
logic [31:0] inst8_p24;
logic [31:0] inst8_p25;
logic [31:0] inst8_p26;
logic [31:0] inst8_p27;
logic [31:0] inst8_p28;
logic [31:0] inst8_p29;
logic [31:0] inst8_p30;
logic [31:0] inst8_p31;
logic [31:0] inst8_p32;
logic [31:0] inst8_p33;
logic inst8_reset;
logic inst8_clk;
logic [1023:0] inst9_in;
logic [1023:0] inst9_out;
logic inst9_clk;
logic inst9_reset;
logic inst9_write_en;
logic [1023:0] inst10_p4;
logic [31:0] inst10_p5;
logic [31:0] inst10_p6;
logic [31:0] inst10_p7;
logic [31:0] inst10_p8;
logic [31:0] inst10_p9;
logic [31:0] inst10_p10;
logic [31:0] inst10_p11;
logic [31:0] inst10_p12;
logic [31:0] inst10_p13;
logic [31:0] inst10_p14;
logic [31:0] inst10_p15;
logic [31:0] inst10_p16;
logic [31:0] inst10_p17;
logic [31:0] inst10_p18;
logic [31:0] inst10_p19;
logic [31:0] inst10_p20;
logic [31:0] inst10_p21;
logic [31:0] inst10_p22;
logic [31:0] inst10_p23;
logic [31:0] inst10_p24;
logic [31:0] inst10_p25;
logic [31:0] inst10_p26;
logic [31:0] inst10_p27;
logic [31:0] inst10_p28;
logic [31:0] inst10_p29;
logic [31:0] inst10_p30;
logic [31:0] inst10_p31;
logic [31:0] inst10_p32;
logic [31:0] inst10_p33;
logic [31:0] inst10_p34;
logic [31:0] inst10_p35;
logic [31:0] inst10_p36;
logic inst10_clk;
logic inst10_reset;
logic [31:0] inst11_p5;
logic [31:0] inst11_p6;
logic [31:0] inst11_p7;
logic [31:0] inst11_p8;
logic [31:0] inst11_p9;
logic [31:0] inst11_p10;
logic [31:0] inst11_p11;
logic [31:0] inst11_p12;
logic [31:0] inst11_p13;
logic [31:0] inst11_p14;
logic [31:0] inst11_p15;
logic [31:0] inst11_p16;
logic [31:0] inst11_p17;
logic [31:0] inst11_p18;
logic [31:0] inst11_p19;
logic [31:0] inst11_p20;
logic [31:0] inst11_p21;
logic [31:0] inst11_p22;
logic [31:0] inst11_p23;
logic [31:0] inst11_p24;
logic [31:0] inst11_p25;
logic [31:0] inst11_p26;
logic [31:0] inst11_p27;
logic [31:0] inst11_p28;
logic [31:0] inst11_p29;
logic [31:0] inst11_p30;
logic [31:0] inst11_p31;
logic [31:0] inst11_p32;
logic [31:0] inst11_p33;
logic [31:0] inst11_p34;
logic [31:0] inst11_p35;
logic [31:0] inst11_p36;
logic [1023:0] inst11_p37;
logic inst11_clk;
logic inst11_reset;
logic [31:0] inst12_p5;
logic [31:0] inst12_p6;
logic [31:0] inst12_p7;
logic [31:0] inst12_p8;
logic [31:0] inst12_p9;
logic [31:0] inst12_p10;
logic [31:0] inst12_p11;
logic [31:0] inst12_p12;
logic [31:0] inst12_p13;
logic [31:0] inst12_p14;
logic [31:0] inst12_p15;
logic [31:0] inst12_p16;
logic [31:0] inst12_p17;
logic [31:0] inst12_p18;
logic [31:0] inst12_p19;
logic [31:0] inst12_p20;
logic [31:0] inst12_p21;
logic [31:0] inst12_p22;
logic [31:0] inst12_p23;
logic [31:0] inst12_p24;
logic [31:0] inst12_p25;
logic [31:0] inst12_p26;
logic [31:0] inst12_p27;
logic [31:0] inst12_p28;
logic [31:0] inst12_p29;
logic [31:0] inst12_p30;
logic [31:0] inst12_p31;
logic [31:0] inst12_p32;
logic [31:0] inst12_p33;
logic [31:0] inst12_p34;
logic [31:0] inst12_p35;
logic [31:0] inst12_p36;
logic [1023:0] inst12_p37;
logic inst12_clk;
logic inst12_reset;
logic [1023:0] inst13_p4;
logic [31:0] inst13_p5;
logic [31:0] inst13_p6;
logic [31:0] inst13_p7;
logic [31:0] inst13_p8;
logic [31:0] inst13_p9;
logic [31:0] inst13_p10;
logic [31:0] inst13_p11;
logic [31:0] inst13_p12;
logic [31:0] inst13_p13;
logic [31:0] inst13_p14;
logic [31:0] inst13_p15;
logic [31:0] inst13_p16;
logic [31:0] inst13_p17;
logic [31:0] inst13_p18;
logic [31:0] inst13_p19;
logic [31:0] inst13_p20;
logic [31:0] inst13_p21;
logic [31:0] inst13_p22;
logic [31:0] inst13_p23;
logic [31:0] inst13_p24;
logic [31:0] inst13_p25;
logic [31:0] inst13_p26;
logic [31:0] inst13_p27;
logic [31:0] inst13_p28;
logic [31:0] inst13_p29;
logic [31:0] inst13_p30;
logic [31:0] inst13_p31;
logic [31:0] inst13_p32;
logic [31:0] inst13_p33;
logic [31:0] inst13_p34;
logic [31:0] inst13_p35;
logic [31:0] inst13_p36;
logic inst13_clk;
logic inst13_reset;
logic [1023:0] inst14_p4;
logic [31:0] inst14_p5;
logic [31:0] inst14_p6;
logic [31:0] inst14_p7;
logic [31:0] inst14_p8;
logic [31:0] inst14_p9;
logic [31:0] inst14_p10;
logic [31:0] inst14_p11;
logic [31:0] inst14_p12;
logic [31:0] inst14_p13;
logic [31:0] inst14_p14;
logic [31:0] inst14_p15;
logic [31:0] inst14_p16;
logic [31:0] inst14_p17;
logic [31:0] inst14_p18;
logic [31:0] inst14_p19;
logic [31:0] inst14_p20;
logic [31:0] inst14_p21;
logic [31:0] inst14_p22;
logic [31:0] inst14_p23;
logic [31:0] inst14_p24;
logic [31:0] inst14_p25;
logic [31:0] inst14_p26;
logic [31:0] inst14_p27;
logic [31:0] inst14_p28;
logic [31:0] inst14_p29;
logic [31:0] inst14_p30;
logic [31:0] inst14_p31;
logic [31:0] inst14_p32;
logic [31:0] inst14_p33;
logic [31:0] inst14_p34;
logic [31:0] inst14_p35;
logic [31:0] inst14_p36;
logic inst14_clk;
logic inst14_reset;
logic [31:0] inst15_p5;
logic [31:0] inst15_p6;
logic [31:0] inst15_p7;
logic [31:0] inst15_p8;
logic [31:0] inst15_p9;
logic [31:0] inst15_p10;
logic [31:0] inst15_p11;
logic [31:0] inst15_p12;
logic [31:0] inst15_p13;
logic [31:0] inst15_p14;
logic [31:0] inst15_p15;
logic [31:0] inst15_p16;
logic [31:0] inst15_p17;
logic [31:0] inst15_p18;
logic [31:0] inst15_p19;
logic [31:0] inst15_p20;
logic [31:0] inst15_p21;
logic [31:0] inst15_p22;
logic [31:0] inst15_p23;
logic [31:0] inst15_p24;
logic [31:0] inst15_p25;
logic [31:0] inst15_p26;
logic [31:0] inst15_p27;
logic [31:0] inst15_p28;
logic [31:0] inst15_p29;
logic [31:0] inst15_p30;
logic [31:0] inst15_p31;
logic [31:0] inst15_p32;
logic [31:0] inst15_p33;
logic [31:0] inst15_p34;
logic [31:0] inst15_p35;
logic [31:0] inst15_p36;
logic [1023:0] inst15_p37;
logic inst15_clk;
logic inst15_reset;
logic [31:0] inst16_p5;
logic [31:0] inst16_p6;
logic [31:0] inst16_p7;
logic [31:0] inst16_p8;
logic [31:0] inst16_p9;
logic [31:0] inst16_p10;
logic [31:0] inst16_p11;
logic [31:0] inst16_p12;
logic [31:0] inst16_p13;
logic [31:0] inst16_p14;
logic [31:0] inst16_p15;
logic [31:0] inst16_p16;
logic [31:0] inst16_p17;
logic [31:0] inst16_p18;
logic [31:0] inst16_p19;
logic [31:0] inst16_p20;
logic [31:0] inst16_p21;
logic [31:0] inst16_p22;
logic [31:0] inst16_p23;
logic [31:0] inst16_p24;
logic [31:0] inst16_p25;
logic [31:0] inst16_p26;
logic [31:0] inst16_p27;
logic [31:0] inst16_p28;
logic [31:0] inst16_p29;
logic [31:0] inst16_p30;
logic [31:0] inst16_p31;
logic [31:0] inst16_p32;
logic [31:0] inst16_p33;
logic [31:0] inst16_p34;
logic [31:0] inst16_p35;
logic [31:0] inst16_p36;
logic [1023:0] inst16_p37;
logic inst16_clk;
logic inst16_reset;
logic [1023:0] inst17_p4;
logic [31:0] inst17_p5;
logic [31:0] inst17_p6;
logic [31:0] inst17_p7;
logic [31:0] inst17_p8;
logic [31:0] inst17_p9;
logic [31:0] inst17_p10;
logic [31:0] inst17_p11;
logic [31:0] inst17_p12;
logic [31:0] inst17_p13;
logic [31:0] inst17_p14;
logic [31:0] inst17_p15;
logic [31:0] inst17_p16;
logic [31:0] inst17_p17;
logic [31:0] inst17_p18;
logic [31:0] inst17_p19;
logic [31:0] inst17_p20;
logic [31:0] inst17_p21;
logic [31:0] inst17_p22;
logic [31:0] inst17_p23;
logic [31:0] inst17_p24;
logic [31:0] inst17_p25;
logic [31:0] inst17_p26;
logic [31:0] inst17_p27;
logic [31:0] inst17_p28;
logic [31:0] inst17_p29;
logic [31:0] inst17_p30;
logic [31:0] inst17_p31;
logic [31:0] inst17_p32;
logic [31:0] inst17_p33;
logic [31:0] inst17_p34;
logic [31:0] inst17_p35;
logic [31:0] inst17_p36;
logic inst17_clk;
logic inst17_reset;
logic [1023:0] inst18_p4;
logic [31:0] inst18_p5;
logic [31:0] inst18_p6;
logic [31:0] inst18_p7;
logic [31:0] inst18_p8;
logic [31:0] inst18_p9;
logic [31:0] inst18_p10;
logic [31:0] inst18_p11;
logic [31:0] inst18_p12;
logic [31:0] inst18_p13;
logic [31:0] inst18_p14;
logic [31:0] inst18_p15;
logic [31:0] inst18_p16;
logic [31:0] inst18_p17;
logic [31:0] inst18_p18;
logic [31:0] inst18_p19;
logic [31:0] inst18_p20;
logic [31:0] inst18_p21;
logic [31:0] inst18_p22;
logic [31:0] inst18_p23;
logic [31:0] inst18_p24;
logic [31:0] inst18_p25;
logic [31:0] inst18_p26;
logic [31:0] inst18_p27;
logic [31:0] inst18_p28;
logic [31:0] inst18_p29;
logic [31:0] inst18_p30;
logic [31:0] inst18_p31;
logic [31:0] inst18_p32;
logic [31:0] inst18_p33;
logic [31:0] inst18_p34;
logic [31:0] inst18_p35;
logic [31:0] inst18_p36;
logic inst18_clk;
logic inst18_reset;
logic [31:0] inst19_p5;
logic [31:0] inst19_p6;
logic [31:0] inst19_p7;
logic [31:0] inst19_p8;
logic [31:0] inst19_p9;
logic [31:0] inst19_p10;
logic [31:0] inst19_p11;
logic [31:0] inst19_p12;
logic [31:0] inst19_p13;
logic [31:0] inst19_p14;
logic [31:0] inst19_p15;
logic [31:0] inst19_p16;
logic [31:0] inst19_p17;
logic [31:0] inst19_p18;
logic [31:0] inst19_p19;
logic [31:0] inst19_p20;
logic [31:0] inst19_p21;
logic [31:0] inst19_p22;
logic [31:0] inst19_p23;
logic [31:0] inst19_p24;
logic [31:0] inst19_p25;
logic [31:0] inst19_p26;
logic [31:0] inst19_p27;
logic [31:0] inst19_p28;
logic [31:0] inst19_p29;
logic [31:0] inst19_p30;
logic [31:0] inst19_p31;
logic [31:0] inst19_p32;
logic [31:0] inst19_p33;
logic [31:0] inst19_p34;
logic [31:0] inst19_p35;
logic [31:0] inst19_p36;
logic [1023:0] inst19_p37;
logic inst19_clk;
logic inst19_reset;
logic [31:0] inst20_p5;
logic [31:0] inst20_p6;
logic [31:0] inst20_p7;
logic [31:0] inst20_p8;
logic [31:0] inst20_p9;
logic [31:0] inst20_p10;
logic [31:0] inst20_p11;
logic [31:0] inst20_p12;
logic [31:0] inst20_p13;
logic [31:0] inst20_p14;
logic [31:0] inst20_p15;
logic [31:0] inst20_p16;
logic [31:0] inst20_p17;
logic [31:0] inst20_p18;
logic [31:0] inst20_p19;
logic [31:0] inst20_p20;
logic [31:0] inst20_p21;
logic [31:0] inst20_p22;
logic [31:0] inst20_p23;
logic [31:0] inst20_p24;
logic [31:0] inst20_p25;
logic [31:0] inst20_p26;
logic [31:0] inst20_p27;
logic [31:0] inst20_p28;
logic [31:0] inst20_p29;
logic [31:0] inst20_p30;
logic [31:0] inst20_p31;
logic [31:0] inst20_p32;
logic [31:0] inst20_p33;
logic [31:0] inst20_p34;
logic [31:0] inst20_p35;
logic [31:0] inst20_p36;
logic [1023:0] inst20_p37;
logic inst20_clk;
logic inst20_reset;
logic [1023:0] inst21_p4;
logic [31:0] inst21_p5;
logic [31:0] inst21_p6;
logic [31:0] inst21_p7;
logic [31:0] inst21_p8;
logic [31:0] inst21_p9;
logic [31:0] inst21_p10;
logic [31:0] inst21_p11;
logic [31:0] inst21_p12;
logic [31:0] inst21_p13;
logic [31:0] inst21_p14;
logic [31:0] inst21_p15;
logic [31:0] inst21_p16;
logic [31:0] inst21_p17;
logic [31:0] inst21_p18;
logic [31:0] inst21_p19;
logic [31:0] inst21_p20;
logic [31:0] inst21_p21;
logic [31:0] inst21_p22;
logic [31:0] inst21_p23;
logic [31:0] inst21_p24;
logic [31:0] inst21_p25;
logic [31:0] inst21_p26;
logic [31:0] inst21_p27;
logic [31:0] inst21_p28;
logic [31:0] inst21_p29;
logic [31:0] inst21_p30;
logic [31:0] inst21_p31;
logic [31:0] inst21_p32;
logic [31:0] inst21_p33;
logic [31:0] inst21_p34;
logic [31:0] inst21_p35;
logic [31:0] inst21_p36;
logic inst21_clk;
logic inst21_reset;
logic [1023:0] inst22_p4;
logic [31:0] inst22_p5;
logic [31:0] inst22_p6;
logic [31:0] inst22_p7;
logic [31:0] inst22_p8;
logic [31:0] inst22_p9;
logic [31:0] inst22_p10;
logic [31:0] inst22_p11;
logic [31:0] inst22_p12;
logic [31:0] inst22_p13;
logic [31:0] inst22_p14;
logic [31:0] inst22_p15;
logic [31:0] inst22_p16;
logic [31:0] inst22_p17;
logic [31:0] inst22_p18;
logic [31:0] inst22_p19;
logic [31:0] inst22_p20;
logic [31:0] inst22_p21;
logic [31:0] inst22_p22;
logic [31:0] inst22_p23;
logic [31:0] inst22_p24;
logic [31:0] inst22_p25;
logic [31:0] inst22_p26;
logic [31:0] inst22_p27;
logic [31:0] inst22_p28;
logic [31:0] inst22_p29;
logic [31:0] inst22_p30;
logic [31:0] inst22_p31;
logic [31:0] inst22_p32;
logic [31:0] inst22_p33;
logic [31:0] inst22_p34;
logic [31:0] inst22_p35;
logic [31:0] inst22_p36;
logic inst22_clk;
logic inst22_reset;
logic [31:0] inst23_p5;
logic [31:0] inst23_p6;
logic [31:0] inst23_p7;
logic [31:0] inst23_p8;
logic [31:0] inst23_p9;
logic [31:0] inst23_p10;
logic [31:0] inst23_p11;
logic [31:0] inst23_p12;
logic [31:0] inst23_p13;
logic [31:0] inst23_p14;
logic [31:0] inst23_p15;
logic [31:0] inst23_p16;
logic [31:0] inst23_p17;
logic [31:0] inst23_p18;
logic [31:0] inst23_p19;
logic [31:0] inst23_p20;
logic [31:0] inst23_p21;
logic [31:0] inst23_p22;
logic [31:0] inst23_p23;
logic [31:0] inst23_p24;
logic [31:0] inst23_p25;
logic [31:0] inst23_p26;
logic [31:0] inst23_p27;
logic [31:0] inst23_p28;
logic [31:0] inst23_p29;
logic [31:0] inst23_p30;
logic [31:0] inst23_p31;
logic [31:0] inst23_p32;
logic [31:0] inst23_p33;
logic [31:0] inst23_p34;
logic [31:0] inst23_p35;
logic [31:0] inst23_p36;
logic [1023:0] inst23_p37;
logic inst23_clk;
logic inst23_reset;
logic [31:0] inst24_p5;
logic [31:0] inst24_p6;
logic [31:0] inst24_p7;
logic [31:0] inst24_p8;
logic [31:0] inst24_p9;
logic [31:0] inst24_p10;
logic [31:0] inst24_p11;
logic [31:0] inst24_p12;
logic [31:0] inst24_p13;
logic [31:0] inst24_p14;
logic [31:0] inst24_p15;
logic [31:0] inst24_p16;
logic [31:0] inst24_p17;
logic [31:0] inst24_p18;
logic [31:0] inst24_p19;
logic [31:0] inst24_p20;
logic [31:0] inst24_p21;
logic [31:0] inst24_p22;
logic [31:0] inst24_p23;
logic [31:0] inst24_p24;
logic [31:0] inst24_p25;
logic [31:0] inst24_p26;
logic [31:0] inst24_p27;
logic [31:0] inst24_p28;
logic [31:0] inst24_p29;
logic [31:0] inst24_p30;
logic [31:0] inst24_p31;
logic [31:0] inst24_p32;
logic [31:0] inst24_p33;
logic [31:0] inst24_p34;
logic [31:0] inst24_p35;
logic [31:0] inst24_p36;
logic [1023:0] inst24_p37;
logic inst24_clk;
logic inst24_reset;
logic [1023:0] inst25_p4;
logic [31:0] inst25_p5;
logic [31:0] inst25_p6;
logic [31:0] inst25_p7;
logic [31:0] inst25_p8;
logic [31:0] inst25_p9;
logic [31:0] inst25_p10;
logic [31:0] inst25_p11;
logic [31:0] inst25_p12;
logic [31:0] inst25_p13;
logic [31:0] inst25_p14;
logic [31:0] inst25_p15;
logic [31:0] inst25_p16;
logic [31:0] inst25_p17;
logic [31:0] inst25_p18;
logic [31:0] inst25_p19;
logic [31:0] inst25_p20;
logic [31:0] inst25_p21;
logic [31:0] inst25_p22;
logic [31:0] inst25_p23;
logic [31:0] inst25_p24;
logic [31:0] inst25_p25;
logic [31:0] inst25_p26;
logic [31:0] inst25_p27;
logic [31:0] inst25_p28;
logic [31:0] inst25_p29;
logic [31:0] inst25_p30;
logic [31:0] inst25_p31;
logic [31:0] inst25_p32;
logic [31:0] inst25_p33;
logic [31:0] inst25_p34;
logic [31:0] inst25_p35;
logic [31:0] inst25_p36;
logic inst25_clk;
logic inst25_reset;
logic [31:0] inst26_p5;
logic [31:0] inst26_p6;
logic [31:0] inst26_p7;
logic [31:0] inst26_p8;
logic [31:0] inst26_p9;
logic [31:0] inst26_p10;
logic [31:0] inst26_p11;
logic [31:0] inst26_p12;
logic [31:0] inst26_p13;
logic [31:0] inst26_p14;
logic [31:0] inst26_p15;
logic [31:0] inst26_p16;
logic [31:0] inst26_p17;
logic [31:0] inst26_p18;
logic [31:0] inst26_p19;
logic [31:0] inst26_p20;
logic [31:0] inst26_p21;
logic [31:0] inst26_p22;
logic [31:0] inst26_p23;
logic [31:0] inst26_p24;
logic [31:0] inst26_p25;
logic [31:0] inst26_p26;
logic [31:0] inst26_p27;
logic [31:0] inst26_p28;
logic [31:0] inst26_p29;
logic [31:0] inst26_p30;
logic [31:0] inst26_p31;
logic [31:0] inst26_p32;
logic [31:0] inst26_p33;
logic [31:0] inst26_p34;
logic [31:0] inst26_p35;
logic [31:0] inst26_p36;
logic [1023:0] inst26_p37;
logic inst26_clk;
logic inst26_reset;
logic [1023:0] inst27_p4;
logic [31:0] inst27_p5;
logic [31:0] inst27_p6;
logic [31:0] inst27_p7;
logic [31:0] inst27_p8;
logic [31:0] inst27_p9;
logic [31:0] inst27_p10;
logic [31:0] inst27_p11;
logic [31:0] inst27_p12;
logic [31:0] inst27_p13;
logic [31:0] inst27_p14;
logic [31:0] inst27_p15;
logic [31:0] inst27_p16;
logic [31:0] inst27_p17;
logic [31:0] inst27_p18;
logic [31:0] inst27_p19;
logic [31:0] inst27_p20;
logic [31:0] inst27_p21;
logic [31:0] inst27_p22;
logic [31:0] inst27_p23;
logic [31:0] inst27_p24;
logic [31:0] inst27_p25;
logic [31:0] inst27_p26;
logic [31:0] inst27_p27;
logic [31:0] inst27_p28;
logic [31:0] inst27_p29;
logic [31:0] inst27_p30;
logic [31:0] inst27_p31;
logic [31:0] inst27_p32;
logic [31:0] inst27_p33;
logic [31:0] inst27_p34;
logic [31:0] inst27_p35;
logic [31:0] inst27_p36;
logic inst27_clk;
logic inst27_reset;
logic [31:0] inst28_p5;
logic [31:0] inst28_p6;
logic [31:0] inst28_p7;
logic [31:0] inst28_p8;
logic [31:0] inst28_p9;
logic [31:0] inst28_p10;
logic [31:0] inst28_p11;
logic [31:0] inst28_p12;
logic [31:0] inst28_p13;
logic [31:0] inst28_p14;
logic [31:0] inst28_p15;
logic [31:0] inst28_p16;
logic [31:0] inst28_p17;
logic [31:0] inst28_p18;
logic [31:0] inst28_p19;
logic [31:0] inst28_p20;
logic [31:0] inst28_p21;
logic [31:0] inst28_p22;
logic [31:0] inst28_p23;
logic [31:0] inst28_p24;
logic [31:0] inst28_p25;
logic [31:0] inst28_p26;
logic [31:0] inst28_p27;
logic [31:0] inst28_p28;
logic [31:0] inst28_p29;
logic [31:0] inst28_p30;
logic [31:0] inst28_p31;
logic [31:0] inst28_p32;
logic [31:0] inst28_p33;
logic [31:0] inst28_p34;
logic [31:0] inst28_p35;
logic [31:0] inst28_p36;
logic [1023:0] inst28_p37;
logic inst28_clk;
logic inst28_reset;
logic [1023:0] inst29_p4;
logic [31:0] inst29_p5;
logic [31:0] inst29_p6;
logic [31:0] inst29_p7;
logic [31:0] inst29_p8;
logic [31:0] inst29_p9;
logic [31:0] inst29_p10;
logic [31:0] inst29_p11;
logic [31:0] inst29_p12;
logic [31:0] inst29_p13;
logic [31:0] inst29_p14;
logic [31:0] inst29_p15;
logic [31:0] inst29_p16;
logic [31:0] inst29_p17;
logic [31:0] inst29_p18;
logic [31:0] inst29_p19;
logic [31:0] inst29_p20;
logic [31:0] inst29_p21;
logic [31:0] inst29_p22;
logic [31:0] inst29_p23;
logic [31:0] inst29_p24;
logic [31:0] inst29_p25;
logic [31:0] inst29_p26;
logic [31:0] inst29_p27;
logic [31:0] inst29_p28;
logic [31:0] inst29_p29;
logic [31:0] inst29_p30;
logic [31:0] inst29_p31;
logic [31:0] inst29_p32;
logic [31:0] inst29_p33;
logic [31:0] inst29_p34;
logic [31:0] inst29_p35;
logic [31:0] inst29_p36;
logic inst29_clk;
logic inst29_reset;
logic [31:0] inst30_p5;
logic [31:0] inst30_p6;
logic [31:0] inst30_p7;
logic [31:0] inst30_p8;
logic [31:0] inst30_p9;
logic [31:0] inst30_p10;
logic [31:0] inst30_p11;
logic [31:0] inst30_p12;
logic [31:0] inst30_p13;
logic [31:0] inst30_p14;
logic [31:0] inst30_p15;
logic [31:0] inst30_p16;
logic [31:0] inst30_p17;
logic [31:0] inst30_p18;
logic [31:0] inst30_p19;
logic [31:0] inst30_p20;
logic [31:0] inst30_p21;
logic [31:0] inst30_p22;
logic [31:0] inst30_p23;
logic [31:0] inst30_p24;
logic [31:0] inst30_p25;
logic [31:0] inst30_p26;
logic [31:0] inst30_p27;
logic [31:0] inst30_p28;
logic [31:0] inst30_p29;
logic [31:0] inst30_p30;
logic [31:0] inst30_p31;
logic [31:0] inst30_p32;
logic [31:0] inst30_p33;
logic [31:0] inst30_p34;
logic [31:0] inst30_p35;
logic [31:0] inst30_p36;
logic [1023:0] inst30_p37;
logic inst30_clk;
logic inst30_reset;
logic [1023:0] inst31_p4;
logic [31:0] inst31_p5;
logic [31:0] inst31_p6;
logic [31:0] inst31_p7;
logic [31:0] inst31_p8;
logic [31:0] inst31_p9;
logic [31:0] inst31_p10;
logic [31:0] inst31_p11;
logic [31:0] inst31_p12;
logic [31:0] inst31_p13;
logic [31:0] inst31_p14;
logic [31:0] inst31_p15;
logic [31:0] inst31_p16;
logic [31:0] inst31_p17;
logic [31:0] inst31_p18;
logic [31:0] inst31_p19;
logic [31:0] inst31_p20;
logic [31:0] inst31_p21;
logic [31:0] inst31_p22;
logic [31:0] inst31_p23;
logic [31:0] inst31_p24;
logic [31:0] inst31_p25;
logic [31:0] inst31_p26;
logic [31:0] inst31_p27;
logic [31:0] inst31_p28;
logic [31:0] inst31_p29;
logic [31:0] inst31_p30;
logic [31:0] inst31_p31;
logic [31:0] inst31_p32;
logic [31:0] inst31_p33;
logic [31:0] inst31_p34;
logic [31:0] inst31_p35;
logic [31:0] inst31_p36;
logic inst31_clk;
logic inst31_reset;
logic [31:0] inst32_p5;
logic [31:0] inst32_p6;
logic [31:0] inst32_p7;
logic [31:0] inst32_p8;
logic [31:0] inst32_p9;
logic [31:0] inst32_p10;
logic [31:0] inst32_p11;
logic [31:0] inst32_p12;
logic [31:0] inst32_p13;
logic [31:0] inst32_p14;
logic [31:0] inst32_p15;
logic [31:0] inst32_p16;
logic [31:0] inst32_p17;
logic [31:0] inst32_p18;
logic [31:0] inst32_p19;
logic [31:0] inst32_p20;
logic [31:0] inst32_p21;
logic [31:0] inst32_p22;
logic [31:0] inst32_p23;
logic [31:0] inst32_p24;
logic [31:0] inst32_p25;
logic [31:0] inst32_p26;
logic [31:0] inst32_p27;
logic [31:0] inst32_p28;
logic [31:0] inst32_p29;
logic [31:0] inst32_p30;
logic [31:0] inst32_p31;
logic [31:0] inst32_p32;
logic [31:0] inst32_p33;
logic [31:0] inst32_p34;
logic [31:0] inst32_p35;
logic [31:0] inst32_p36;
logic [1023:0] inst32_p37;
logic inst32_clk;
logic inst32_reset;
logic [1023:0] inst33_p4;
logic [31:0] inst33_p5;
logic [31:0] inst33_p6;
logic [31:0] inst33_p7;
logic [31:0] inst33_p8;
logic [31:0] inst33_p9;
logic [31:0] inst33_p10;
logic [31:0] inst33_p11;
logic [31:0] inst33_p12;
logic [31:0] inst33_p13;
logic [31:0] inst33_p14;
logic [31:0] inst33_p15;
logic [31:0] inst33_p16;
logic [31:0] inst33_p17;
logic [31:0] inst33_p18;
logic [31:0] inst33_p19;
logic [31:0] inst33_p20;
logic [31:0] inst33_p21;
logic [31:0] inst33_p22;
logic [31:0] inst33_p23;
logic [31:0] inst33_p24;
logic [31:0] inst33_p25;
logic [31:0] inst33_p26;
logic [31:0] inst33_p27;
logic [31:0] inst33_p28;
logic [31:0] inst33_p29;
logic [31:0] inst33_p30;
logic [31:0] inst33_p31;
logic [31:0] inst33_p32;
logic [31:0] inst33_p33;
logic [31:0] inst33_p34;
logic [31:0] inst33_p35;
logic [31:0] inst33_p36;
logic inst33_clk;
logic inst33_reset;
counter_chain_2_128 ev00 (
    ._0_0(ev00__0_0),
    ._0state(ev00__0state),
    ._1_0(ev00__1_0),
    ._1state(ev00__1state),
    .clk(ev00_clk),
    .done(ev00_done),
    .go(ev00_go),
    .reset(ev00_reset)
);
comp35 inst0 (
    .clk(inst0_clk),
    .ev0(inst0_ev0),
    .p100(inst0_p100),
    .p101(inst0_p101),
    .p102(inst0_p102),
    .p103(inst0_p103),
    .p104(inst0_p104),
    .p105(inst0_p105),
    .p106(inst0_p106),
    .p107(inst0_p107),
    .p108(inst0_p108),
    .p109(inst0_p109),
    .p110(inst0_p110),
    .p111(inst0_p111),
    .p112(inst0_p112),
    .p113(inst0_p113),
    .p114(inst0_p114),
    .p115(inst0_p115),
    .p116(inst0_p116),
    .p117(inst0_p117),
    .p118(inst0_p118),
    .p119(inst0_p119),
    .p120(inst0_p120),
    .p121(inst0_p121),
    .p122(inst0_p122),
    .p43(inst0_p43),
    .p44(inst0_p44),
    .p45(inst0_p45),
    .p46(inst0_p46),
    .p47(inst0_p47),
    .p48(inst0_p48),
    .p49(inst0_p49),
    .p50(inst0_p50),
    .p51(inst0_p51),
    .p52(inst0_p52),
    .p53(inst0_p53),
    .p54(inst0_p54),
    .p55(inst0_p55),
    .p56(inst0_p56),
    .p57(inst0_p57),
    .p58(inst0_p58),
    .p59(inst0_p59),
    .p60(inst0_p60),
    .p61(inst0_p61),
    .p62(inst0_p62),
    .p63(inst0_p63),
    .p64(inst0_p64),
    .p65(inst0_p65),
    .p66(inst0_p66),
    .p67(inst0_p67),
    .p68(inst0_p68),
    .p69(inst0_p69),
    .p70(inst0_p70),
    .p71(inst0_p71),
    .p72(inst0_p72),
    .p73(inst0_p73),
    .p74(inst0_p74),
    .p75(inst0_p75),
    .p76(inst0_p76),
    .p77(inst0_p77),
    .p78(inst0_p78),
    .p79(inst0_p79),
    .p80(inst0_p80),
    .p81(inst0_p81),
    .p82(inst0_p82),
    .p83(inst0_p83),
    .p84(inst0_p84),
    .p85(inst0_p85),
    .p86(inst0_p86),
    .p87(inst0_p87),
    .p88(inst0_p88),
    .p89(inst0_p89),
    .p90(inst0_p90),
    .p91(inst0_p91),
    .p92(inst0_p92),
    .p93(inst0_p93),
    .p94(inst0_p94),
    .p95(inst0_p95),
    .p96(inst0_p96),
    .p97(inst0_p97),
    .p98(inst0_p98),
    .p99(inst0_p99),
    .reset(inst0_reset)
);
comp36 inst1 (
    .clk(inst1_clk),
    .p10(inst1_p10),
    .p11(inst1_p11),
    .p12(inst1_p12),
    .p13(inst1_p13),
    .p14(inst1_p14),
    .p15(inst1_p15),
    .p16(inst1_p16),
    .p17(inst1_p17),
    .p18(inst1_p18),
    .p19(inst1_p19),
    .p2(inst1_p2),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .p3(inst1_p3),
    .p30(inst1_p30),
    .p31(inst1_p31),
    .p32(inst1_p32),
    .p33(inst1_p33),
    .p34(inst1_p34),
    .p35(inst1_p35),
    .p36(inst1_p36),
    .p37(inst1_p37),
    .p38(inst1_p38),
    .p39(inst1_p39),
    .p4(inst1_p4),
    .p40(inst1_p40),
    .p41(inst1_p41),
    .p42(inst1_p42),
    .p43(inst1_p43),
    .p44(inst1_p44),
    .p45(inst1_p45),
    .p46(inst1_p46),
    .p47(inst1_p47),
    .p48(inst1_p48),
    .p49(inst1_p49),
    .p5(inst1_p5),
    .p50(inst1_p50),
    .p51(inst1_p51),
    .p52(inst1_p52),
    .p53(inst1_p53),
    .p54(inst1_p54),
    .p55(inst1_p55),
    .p56(inst1_p56),
    .p57(inst1_p57),
    .p58(inst1_p58),
    .p59(inst1_p59),
    .p6(inst1_p6),
    .p60(inst1_p60),
    .p61(inst1_p61),
    .p62(inst1_p62),
    .p63(inst1_p63),
    .p64(inst1_p64),
    .p65(inst1_p65),
    .p7(inst1_p7),
    .p8(inst1_p8),
    .p9(inst1_p9),
    .reset(inst1_reset)
);
comp49 inst2 (
    .clk(inst2_clk),
    .p17(inst2_p17),
    .p18(inst2_p18),
    .p19(inst2_p19),
    .p20(inst2_p20),
    .p21(inst2_p21),
    .p22(inst2_p22),
    .p23(inst2_p23),
    .p24(inst2_p24),
    .p25(inst2_p25),
    .p26(inst2_p26),
    .p27(inst2_p27),
    .p28(inst2_p28),
    .p29(inst2_p29),
    .p30(inst2_p30),
    .p31(inst2_p31),
    .p32(inst2_p32),
    .reset(inst2_reset)
);
comp50 inst3 (
    .clk(inst3_clk),
    .p10(inst3_p10),
    .p11(inst3_p11),
    .p12(inst3_p12),
    .p13(inst3_p13),
    .p14(inst3_p14),
    .p15(inst3_p15),
    .p16(inst3_p16),
    .p17(inst3_p17),
    .p18(inst3_p18),
    .p19(inst3_p19),
    .p2(inst3_p2),
    .p20(inst3_p20),
    .p21(inst3_p21),
    .p22(inst3_p22),
    .p23(inst3_p23),
    .p24(inst3_p24),
    .p25(inst3_p25),
    .p26(inst3_p26),
    .p27(inst3_p27),
    .p28(inst3_p28),
    .p29(inst3_p29),
    .p3(inst3_p3),
    .p30(inst3_p30),
    .p31(inst3_p31),
    .p32(inst3_p32),
    .p33(inst3_p33),
    .p34(inst3_p34),
    .p35(inst3_p35),
    .p36(inst3_p36),
    .p37(inst3_p37),
    .p38(inst3_p38),
    .p39(inst3_p39),
    .p4(inst3_p4),
    .p40(inst3_p40),
    .p41(inst3_p41),
    .p42(inst3_p42),
    .p43(inst3_p43),
    .p44(inst3_p44),
    .p45(inst3_p45),
    .p46(inst3_p46),
    .p47(inst3_p47),
    .p48(inst3_p48),
    .p49(inst3_p49),
    .p5(inst3_p5),
    .p50(inst3_p50),
    .p51(inst3_p51),
    .p52(inst3_p52),
    .p53(inst3_p53),
    .p54(inst3_p54),
    .p55(inst3_p55),
    .p56(inst3_p56),
    .p57(inst3_p57),
    .p58(inst3_p58),
    .p59(inst3_p59),
    .p6(inst3_p6),
    .p60(inst3_p60),
    .p61(inst3_p61),
    .p62(inst3_p62),
    .p63(inst3_p63),
    .p64(inst3_p64),
    .p65(inst3_p65),
    .p7(inst3_p7),
    .p8(inst3_p8),
    .p9(inst3_p9),
    .reset(inst3_reset)
);
Delay # (
    .WIDTH(1024)
) inst4 (
    .clk(inst4_clk),
    .in(inst4_in),
    .out(inst4_out),
    .reset(inst4_reset)
);
comp52 inst5 (
    .clk(inst5_clk),
    .p10(inst5_p10),
    .p11(inst5_p11),
    .p12(inst5_p12),
    .p13(inst5_p13),
    .p14(inst5_p14),
    .p15(inst5_p15),
    .p16(inst5_p16),
    .p17(inst5_p17),
    .p18(inst5_p18),
    .p19(inst5_p19),
    .p2(inst5_p2),
    .p20(inst5_p20),
    .p21(inst5_p21),
    .p22(inst5_p22),
    .p23(inst5_p23),
    .p24(inst5_p24),
    .p25(inst5_p25),
    .p26(inst5_p26),
    .p27(inst5_p27),
    .p28(inst5_p28),
    .p29(inst5_p29),
    .p3(inst5_p3),
    .p30(inst5_p30),
    .p31(inst5_p31),
    .p32(inst5_p32),
    .p33(inst5_p33),
    .p4(inst5_p4),
    .p5(inst5_p5),
    .p6(inst5_p6),
    .p7(inst5_p7),
    .p8(inst5_p8),
    .p9(inst5_p9),
    .reset(inst5_reset)
);
comp53 inst6 (
    .clk(inst6_clk),
    .p10(inst6_p10),
    .p11(inst6_p11),
    .p12(inst6_p12),
    .p13(inst6_p13),
    .p14(inst6_p14),
    .p15(inst6_p15),
    .p16(inst6_p16),
    .p17(inst6_p17),
    .p18(inst6_p18),
    .p19(inst6_p19),
    .p2(inst6_p2),
    .p20(inst6_p20),
    .p21(inst6_p21),
    .p22(inst6_p22),
    .p23(inst6_p23),
    .p24(inst6_p24),
    .p25(inst6_p25),
    .p26(inst6_p26),
    .p27(inst6_p27),
    .p28(inst6_p28),
    .p29(inst6_p29),
    .p3(inst6_p3),
    .p30(inst6_p30),
    .p31(inst6_p31),
    .p32(inst6_p32),
    .p33(inst6_p33),
    .p4(inst6_p4),
    .p5(inst6_p5),
    .p6(inst6_p6),
    .p7(inst6_p7),
    .p8(inst6_p8),
    .p9(inst6_p9),
    .reset(inst6_reset)
);
comp54 inst7 (
    .clk(inst7_clk),
    .p10(inst7_p10),
    .p11(inst7_p11),
    .p12(inst7_p12),
    .p13(inst7_p13),
    .p14(inst7_p14),
    .p15(inst7_p15),
    .p16(inst7_p16),
    .p17(inst7_p17),
    .p18(inst7_p18),
    .p19(inst7_p19),
    .p2(inst7_p2),
    .p20(inst7_p20),
    .p21(inst7_p21),
    .p22(inst7_p22),
    .p23(inst7_p23),
    .p24(inst7_p24),
    .p25(inst7_p25),
    .p26(inst7_p26),
    .p27(inst7_p27),
    .p28(inst7_p28),
    .p29(inst7_p29),
    .p3(inst7_p3),
    .p30(inst7_p30),
    .p31(inst7_p31),
    .p32(inst7_p32),
    .p33(inst7_p33),
    .p4(inst7_p4),
    .p5(inst7_p5),
    .p6(inst7_p6),
    .p7(inst7_p7),
    .p8(inst7_p8),
    .p9(inst7_p9),
    .reset(inst7_reset)
);
comp55 inst8 (
    .clk(inst8_clk),
    .p10(inst8_p10),
    .p11(inst8_p11),
    .p12(inst8_p12),
    .p13(inst8_p13),
    .p14(inst8_p14),
    .p15(inst8_p15),
    .p16(inst8_p16),
    .p17(inst8_p17),
    .p18(inst8_p18),
    .p19(inst8_p19),
    .p2(inst8_p2),
    .p20(inst8_p20),
    .p21(inst8_p21),
    .p22(inst8_p22),
    .p23(inst8_p23),
    .p24(inst8_p24),
    .p25(inst8_p25),
    .p26(inst8_p26),
    .p27(inst8_p27),
    .p28(inst8_p28),
    .p29(inst8_p29),
    .p3(inst8_p3),
    .p30(inst8_p30),
    .p31(inst8_p31),
    .p32(inst8_p32),
    .p33(inst8_p33),
    .p4(inst8_p4),
    .p5(inst8_p5),
    .p6(inst8_p6),
    .p7(inst8_p7),
    .p8(inst8_p8),
    .p9(inst8_p9),
    .reset(inst8_reset)
);
PassThroughRegister # (
    .WIDTH(1024)
) inst9 (
    .clk(inst9_clk),
    .in(inst9_in),
    .out(inst9_out),
    .reset(inst9_reset),
    .write_en(inst9_write_en)
);
comp57 inst10 (
    .clk(inst10_clk),
    .p10(inst10_p10),
    .p11(inst10_p11),
    .p12(inst10_p12),
    .p13(inst10_p13),
    .p14(inst10_p14),
    .p15(inst10_p15),
    .p16(inst10_p16),
    .p17(inst10_p17),
    .p18(inst10_p18),
    .p19(inst10_p19),
    .p20(inst10_p20),
    .p21(inst10_p21),
    .p22(inst10_p22),
    .p23(inst10_p23),
    .p24(inst10_p24),
    .p25(inst10_p25),
    .p26(inst10_p26),
    .p27(inst10_p27),
    .p28(inst10_p28),
    .p29(inst10_p29),
    .p30(inst10_p30),
    .p31(inst10_p31),
    .p32(inst10_p32),
    .p33(inst10_p33),
    .p34(inst10_p34),
    .p35(inst10_p35),
    .p36(inst10_p36),
    .p4(inst10_p4),
    .p5(inst10_p5),
    .p6(inst10_p6),
    .p7(inst10_p7),
    .p8(inst10_p8),
    .p9(inst10_p9),
    .reset(inst10_reset)
);
comp91 inst11 (
    .clk(inst11_clk),
    .p10(inst11_p10),
    .p11(inst11_p11),
    .p12(inst11_p12),
    .p13(inst11_p13),
    .p14(inst11_p14),
    .p15(inst11_p15),
    .p16(inst11_p16),
    .p17(inst11_p17),
    .p18(inst11_p18),
    .p19(inst11_p19),
    .p20(inst11_p20),
    .p21(inst11_p21),
    .p22(inst11_p22),
    .p23(inst11_p23),
    .p24(inst11_p24),
    .p25(inst11_p25),
    .p26(inst11_p26),
    .p27(inst11_p27),
    .p28(inst11_p28),
    .p29(inst11_p29),
    .p30(inst11_p30),
    .p31(inst11_p31),
    .p32(inst11_p32),
    .p33(inst11_p33),
    .p34(inst11_p34),
    .p35(inst11_p35),
    .p36(inst11_p36),
    .p37(inst11_p37),
    .p5(inst11_p5),
    .p6(inst11_p6),
    .p7(inst11_p7),
    .p8(inst11_p8),
    .p9(inst11_p9),
    .reset(inst11_reset)
);
comp91 inst12 (
    .clk(inst12_clk),
    .p10(inst12_p10),
    .p11(inst12_p11),
    .p12(inst12_p12),
    .p13(inst12_p13),
    .p14(inst12_p14),
    .p15(inst12_p15),
    .p16(inst12_p16),
    .p17(inst12_p17),
    .p18(inst12_p18),
    .p19(inst12_p19),
    .p20(inst12_p20),
    .p21(inst12_p21),
    .p22(inst12_p22),
    .p23(inst12_p23),
    .p24(inst12_p24),
    .p25(inst12_p25),
    .p26(inst12_p26),
    .p27(inst12_p27),
    .p28(inst12_p28),
    .p29(inst12_p29),
    .p30(inst12_p30),
    .p31(inst12_p31),
    .p32(inst12_p32),
    .p33(inst12_p33),
    .p34(inst12_p34),
    .p35(inst12_p35),
    .p36(inst12_p36),
    .p37(inst12_p37),
    .p5(inst12_p5),
    .p6(inst12_p6),
    .p7(inst12_p7),
    .p8(inst12_p8),
    .p9(inst12_p9),
    .reset(inst12_reset)
);
comp57 inst13 (
    .clk(inst13_clk),
    .p10(inst13_p10),
    .p11(inst13_p11),
    .p12(inst13_p12),
    .p13(inst13_p13),
    .p14(inst13_p14),
    .p15(inst13_p15),
    .p16(inst13_p16),
    .p17(inst13_p17),
    .p18(inst13_p18),
    .p19(inst13_p19),
    .p20(inst13_p20),
    .p21(inst13_p21),
    .p22(inst13_p22),
    .p23(inst13_p23),
    .p24(inst13_p24),
    .p25(inst13_p25),
    .p26(inst13_p26),
    .p27(inst13_p27),
    .p28(inst13_p28),
    .p29(inst13_p29),
    .p30(inst13_p30),
    .p31(inst13_p31),
    .p32(inst13_p32),
    .p33(inst13_p33),
    .p34(inst13_p34),
    .p35(inst13_p35),
    .p36(inst13_p36),
    .p4(inst13_p4),
    .p5(inst13_p5),
    .p6(inst13_p6),
    .p7(inst13_p7),
    .p8(inst13_p8),
    .p9(inst13_p9),
    .reset(inst13_reset)
);
comp57 inst14 (
    .clk(inst14_clk),
    .p10(inst14_p10),
    .p11(inst14_p11),
    .p12(inst14_p12),
    .p13(inst14_p13),
    .p14(inst14_p14),
    .p15(inst14_p15),
    .p16(inst14_p16),
    .p17(inst14_p17),
    .p18(inst14_p18),
    .p19(inst14_p19),
    .p20(inst14_p20),
    .p21(inst14_p21),
    .p22(inst14_p22),
    .p23(inst14_p23),
    .p24(inst14_p24),
    .p25(inst14_p25),
    .p26(inst14_p26),
    .p27(inst14_p27),
    .p28(inst14_p28),
    .p29(inst14_p29),
    .p30(inst14_p30),
    .p31(inst14_p31),
    .p32(inst14_p32),
    .p33(inst14_p33),
    .p34(inst14_p34),
    .p35(inst14_p35),
    .p36(inst14_p36),
    .p4(inst14_p4),
    .p5(inst14_p5),
    .p6(inst14_p6),
    .p7(inst14_p7),
    .p8(inst14_p8),
    .p9(inst14_p9),
    .reset(inst14_reset)
);
comp91 inst15 (
    .clk(inst15_clk),
    .p10(inst15_p10),
    .p11(inst15_p11),
    .p12(inst15_p12),
    .p13(inst15_p13),
    .p14(inst15_p14),
    .p15(inst15_p15),
    .p16(inst15_p16),
    .p17(inst15_p17),
    .p18(inst15_p18),
    .p19(inst15_p19),
    .p20(inst15_p20),
    .p21(inst15_p21),
    .p22(inst15_p22),
    .p23(inst15_p23),
    .p24(inst15_p24),
    .p25(inst15_p25),
    .p26(inst15_p26),
    .p27(inst15_p27),
    .p28(inst15_p28),
    .p29(inst15_p29),
    .p30(inst15_p30),
    .p31(inst15_p31),
    .p32(inst15_p32),
    .p33(inst15_p33),
    .p34(inst15_p34),
    .p35(inst15_p35),
    .p36(inst15_p36),
    .p37(inst15_p37),
    .p5(inst15_p5),
    .p6(inst15_p6),
    .p7(inst15_p7),
    .p8(inst15_p8),
    .p9(inst15_p9),
    .reset(inst15_reset)
);
comp91 inst16 (
    .clk(inst16_clk),
    .p10(inst16_p10),
    .p11(inst16_p11),
    .p12(inst16_p12),
    .p13(inst16_p13),
    .p14(inst16_p14),
    .p15(inst16_p15),
    .p16(inst16_p16),
    .p17(inst16_p17),
    .p18(inst16_p18),
    .p19(inst16_p19),
    .p20(inst16_p20),
    .p21(inst16_p21),
    .p22(inst16_p22),
    .p23(inst16_p23),
    .p24(inst16_p24),
    .p25(inst16_p25),
    .p26(inst16_p26),
    .p27(inst16_p27),
    .p28(inst16_p28),
    .p29(inst16_p29),
    .p30(inst16_p30),
    .p31(inst16_p31),
    .p32(inst16_p32),
    .p33(inst16_p33),
    .p34(inst16_p34),
    .p35(inst16_p35),
    .p36(inst16_p36),
    .p37(inst16_p37),
    .p5(inst16_p5),
    .p6(inst16_p6),
    .p7(inst16_p7),
    .p8(inst16_p8),
    .p9(inst16_p9),
    .reset(inst16_reset)
);
comp57 inst17 (
    .clk(inst17_clk),
    .p10(inst17_p10),
    .p11(inst17_p11),
    .p12(inst17_p12),
    .p13(inst17_p13),
    .p14(inst17_p14),
    .p15(inst17_p15),
    .p16(inst17_p16),
    .p17(inst17_p17),
    .p18(inst17_p18),
    .p19(inst17_p19),
    .p20(inst17_p20),
    .p21(inst17_p21),
    .p22(inst17_p22),
    .p23(inst17_p23),
    .p24(inst17_p24),
    .p25(inst17_p25),
    .p26(inst17_p26),
    .p27(inst17_p27),
    .p28(inst17_p28),
    .p29(inst17_p29),
    .p30(inst17_p30),
    .p31(inst17_p31),
    .p32(inst17_p32),
    .p33(inst17_p33),
    .p34(inst17_p34),
    .p35(inst17_p35),
    .p36(inst17_p36),
    .p4(inst17_p4),
    .p5(inst17_p5),
    .p6(inst17_p6),
    .p7(inst17_p7),
    .p8(inst17_p8),
    .p9(inst17_p9),
    .reset(inst17_reset)
);
comp57 inst18 (
    .clk(inst18_clk),
    .p10(inst18_p10),
    .p11(inst18_p11),
    .p12(inst18_p12),
    .p13(inst18_p13),
    .p14(inst18_p14),
    .p15(inst18_p15),
    .p16(inst18_p16),
    .p17(inst18_p17),
    .p18(inst18_p18),
    .p19(inst18_p19),
    .p20(inst18_p20),
    .p21(inst18_p21),
    .p22(inst18_p22),
    .p23(inst18_p23),
    .p24(inst18_p24),
    .p25(inst18_p25),
    .p26(inst18_p26),
    .p27(inst18_p27),
    .p28(inst18_p28),
    .p29(inst18_p29),
    .p30(inst18_p30),
    .p31(inst18_p31),
    .p32(inst18_p32),
    .p33(inst18_p33),
    .p34(inst18_p34),
    .p35(inst18_p35),
    .p36(inst18_p36),
    .p4(inst18_p4),
    .p5(inst18_p5),
    .p6(inst18_p6),
    .p7(inst18_p7),
    .p8(inst18_p8),
    .p9(inst18_p9),
    .reset(inst18_reset)
);
comp91 inst19 (
    .clk(inst19_clk),
    .p10(inst19_p10),
    .p11(inst19_p11),
    .p12(inst19_p12),
    .p13(inst19_p13),
    .p14(inst19_p14),
    .p15(inst19_p15),
    .p16(inst19_p16),
    .p17(inst19_p17),
    .p18(inst19_p18),
    .p19(inst19_p19),
    .p20(inst19_p20),
    .p21(inst19_p21),
    .p22(inst19_p22),
    .p23(inst19_p23),
    .p24(inst19_p24),
    .p25(inst19_p25),
    .p26(inst19_p26),
    .p27(inst19_p27),
    .p28(inst19_p28),
    .p29(inst19_p29),
    .p30(inst19_p30),
    .p31(inst19_p31),
    .p32(inst19_p32),
    .p33(inst19_p33),
    .p34(inst19_p34),
    .p35(inst19_p35),
    .p36(inst19_p36),
    .p37(inst19_p37),
    .p5(inst19_p5),
    .p6(inst19_p6),
    .p7(inst19_p7),
    .p8(inst19_p8),
    .p9(inst19_p9),
    .reset(inst19_reset)
);
comp91 inst20 (
    .clk(inst20_clk),
    .p10(inst20_p10),
    .p11(inst20_p11),
    .p12(inst20_p12),
    .p13(inst20_p13),
    .p14(inst20_p14),
    .p15(inst20_p15),
    .p16(inst20_p16),
    .p17(inst20_p17),
    .p18(inst20_p18),
    .p19(inst20_p19),
    .p20(inst20_p20),
    .p21(inst20_p21),
    .p22(inst20_p22),
    .p23(inst20_p23),
    .p24(inst20_p24),
    .p25(inst20_p25),
    .p26(inst20_p26),
    .p27(inst20_p27),
    .p28(inst20_p28),
    .p29(inst20_p29),
    .p30(inst20_p30),
    .p31(inst20_p31),
    .p32(inst20_p32),
    .p33(inst20_p33),
    .p34(inst20_p34),
    .p35(inst20_p35),
    .p36(inst20_p36),
    .p37(inst20_p37),
    .p5(inst20_p5),
    .p6(inst20_p6),
    .p7(inst20_p7),
    .p8(inst20_p8),
    .p9(inst20_p9),
    .reset(inst20_reset)
);
comp57 inst21 (
    .clk(inst21_clk),
    .p10(inst21_p10),
    .p11(inst21_p11),
    .p12(inst21_p12),
    .p13(inst21_p13),
    .p14(inst21_p14),
    .p15(inst21_p15),
    .p16(inst21_p16),
    .p17(inst21_p17),
    .p18(inst21_p18),
    .p19(inst21_p19),
    .p20(inst21_p20),
    .p21(inst21_p21),
    .p22(inst21_p22),
    .p23(inst21_p23),
    .p24(inst21_p24),
    .p25(inst21_p25),
    .p26(inst21_p26),
    .p27(inst21_p27),
    .p28(inst21_p28),
    .p29(inst21_p29),
    .p30(inst21_p30),
    .p31(inst21_p31),
    .p32(inst21_p32),
    .p33(inst21_p33),
    .p34(inst21_p34),
    .p35(inst21_p35),
    .p36(inst21_p36),
    .p4(inst21_p4),
    .p5(inst21_p5),
    .p6(inst21_p6),
    .p7(inst21_p7),
    .p8(inst21_p8),
    .p9(inst21_p9),
    .reset(inst21_reset)
);
comp57 inst22 (
    .clk(inst22_clk),
    .p10(inst22_p10),
    .p11(inst22_p11),
    .p12(inst22_p12),
    .p13(inst22_p13),
    .p14(inst22_p14),
    .p15(inst22_p15),
    .p16(inst22_p16),
    .p17(inst22_p17),
    .p18(inst22_p18),
    .p19(inst22_p19),
    .p20(inst22_p20),
    .p21(inst22_p21),
    .p22(inst22_p22),
    .p23(inst22_p23),
    .p24(inst22_p24),
    .p25(inst22_p25),
    .p26(inst22_p26),
    .p27(inst22_p27),
    .p28(inst22_p28),
    .p29(inst22_p29),
    .p30(inst22_p30),
    .p31(inst22_p31),
    .p32(inst22_p32),
    .p33(inst22_p33),
    .p34(inst22_p34),
    .p35(inst22_p35),
    .p36(inst22_p36),
    .p4(inst22_p4),
    .p5(inst22_p5),
    .p6(inst22_p6),
    .p7(inst22_p7),
    .p8(inst22_p8),
    .p9(inst22_p9),
    .reset(inst22_reset)
);
comp91 inst23 (
    .clk(inst23_clk),
    .p10(inst23_p10),
    .p11(inst23_p11),
    .p12(inst23_p12),
    .p13(inst23_p13),
    .p14(inst23_p14),
    .p15(inst23_p15),
    .p16(inst23_p16),
    .p17(inst23_p17),
    .p18(inst23_p18),
    .p19(inst23_p19),
    .p20(inst23_p20),
    .p21(inst23_p21),
    .p22(inst23_p22),
    .p23(inst23_p23),
    .p24(inst23_p24),
    .p25(inst23_p25),
    .p26(inst23_p26),
    .p27(inst23_p27),
    .p28(inst23_p28),
    .p29(inst23_p29),
    .p30(inst23_p30),
    .p31(inst23_p31),
    .p32(inst23_p32),
    .p33(inst23_p33),
    .p34(inst23_p34),
    .p35(inst23_p35),
    .p36(inst23_p36),
    .p37(inst23_p37),
    .p5(inst23_p5),
    .p6(inst23_p6),
    .p7(inst23_p7),
    .p8(inst23_p8),
    .p9(inst23_p9),
    .reset(inst23_reset)
);
comp91 inst24 (
    .clk(inst24_clk),
    .p10(inst24_p10),
    .p11(inst24_p11),
    .p12(inst24_p12),
    .p13(inst24_p13),
    .p14(inst24_p14),
    .p15(inst24_p15),
    .p16(inst24_p16),
    .p17(inst24_p17),
    .p18(inst24_p18),
    .p19(inst24_p19),
    .p20(inst24_p20),
    .p21(inst24_p21),
    .p22(inst24_p22),
    .p23(inst24_p23),
    .p24(inst24_p24),
    .p25(inst24_p25),
    .p26(inst24_p26),
    .p27(inst24_p27),
    .p28(inst24_p28),
    .p29(inst24_p29),
    .p30(inst24_p30),
    .p31(inst24_p31),
    .p32(inst24_p32),
    .p33(inst24_p33),
    .p34(inst24_p34),
    .p35(inst24_p35),
    .p36(inst24_p36),
    .p37(inst24_p37),
    .p5(inst24_p5),
    .p6(inst24_p6),
    .p7(inst24_p7),
    .p8(inst24_p8),
    .p9(inst24_p9),
    .reset(inst24_reset)
);
comp57 inst25 (
    .clk(inst25_clk),
    .p10(inst25_p10),
    .p11(inst25_p11),
    .p12(inst25_p12),
    .p13(inst25_p13),
    .p14(inst25_p14),
    .p15(inst25_p15),
    .p16(inst25_p16),
    .p17(inst25_p17),
    .p18(inst25_p18),
    .p19(inst25_p19),
    .p20(inst25_p20),
    .p21(inst25_p21),
    .p22(inst25_p22),
    .p23(inst25_p23),
    .p24(inst25_p24),
    .p25(inst25_p25),
    .p26(inst25_p26),
    .p27(inst25_p27),
    .p28(inst25_p28),
    .p29(inst25_p29),
    .p30(inst25_p30),
    .p31(inst25_p31),
    .p32(inst25_p32),
    .p33(inst25_p33),
    .p34(inst25_p34),
    .p35(inst25_p35),
    .p36(inst25_p36),
    .p4(inst25_p4),
    .p5(inst25_p5),
    .p6(inst25_p6),
    .p7(inst25_p7),
    .p8(inst25_p8),
    .p9(inst25_p9),
    .reset(inst25_reset)
);
comp91 inst26 (
    .clk(inst26_clk),
    .p10(inst26_p10),
    .p11(inst26_p11),
    .p12(inst26_p12),
    .p13(inst26_p13),
    .p14(inst26_p14),
    .p15(inst26_p15),
    .p16(inst26_p16),
    .p17(inst26_p17),
    .p18(inst26_p18),
    .p19(inst26_p19),
    .p20(inst26_p20),
    .p21(inst26_p21),
    .p22(inst26_p22),
    .p23(inst26_p23),
    .p24(inst26_p24),
    .p25(inst26_p25),
    .p26(inst26_p26),
    .p27(inst26_p27),
    .p28(inst26_p28),
    .p29(inst26_p29),
    .p30(inst26_p30),
    .p31(inst26_p31),
    .p32(inst26_p32),
    .p33(inst26_p33),
    .p34(inst26_p34),
    .p35(inst26_p35),
    .p36(inst26_p36),
    .p37(inst26_p37),
    .p5(inst26_p5),
    .p6(inst26_p6),
    .p7(inst26_p7),
    .p8(inst26_p8),
    .p9(inst26_p9),
    .reset(inst26_reset)
);
comp57 inst27 (
    .clk(inst27_clk),
    .p10(inst27_p10),
    .p11(inst27_p11),
    .p12(inst27_p12),
    .p13(inst27_p13),
    .p14(inst27_p14),
    .p15(inst27_p15),
    .p16(inst27_p16),
    .p17(inst27_p17),
    .p18(inst27_p18),
    .p19(inst27_p19),
    .p20(inst27_p20),
    .p21(inst27_p21),
    .p22(inst27_p22),
    .p23(inst27_p23),
    .p24(inst27_p24),
    .p25(inst27_p25),
    .p26(inst27_p26),
    .p27(inst27_p27),
    .p28(inst27_p28),
    .p29(inst27_p29),
    .p30(inst27_p30),
    .p31(inst27_p31),
    .p32(inst27_p32),
    .p33(inst27_p33),
    .p34(inst27_p34),
    .p35(inst27_p35),
    .p36(inst27_p36),
    .p4(inst27_p4),
    .p5(inst27_p5),
    .p6(inst27_p6),
    .p7(inst27_p7),
    .p8(inst27_p8),
    .p9(inst27_p9),
    .reset(inst27_reset)
);
comp91 inst28 (
    .clk(inst28_clk),
    .p10(inst28_p10),
    .p11(inst28_p11),
    .p12(inst28_p12),
    .p13(inst28_p13),
    .p14(inst28_p14),
    .p15(inst28_p15),
    .p16(inst28_p16),
    .p17(inst28_p17),
    .p18(inst28_p18),
    .p19(inst28_p19),
    .p20(inst28_p20),
    .p21(inst28_p21),
    .p22(inst28_p22),
    .p23(inst28_p23),
    .p24(inst28_p24),
    .p25(inst28_p25),
    .p26(inst28_p26),
    .p27(inst28_p27),
    .p28(inst28_p28),
    .p29(inst28_p29),
    .p30(inst28_p30),
    .p31(inst28_p31),
    .p32(inst28_p32),
    .p33(inst28_p33),
    .p34(inst28_p34),
    .p35(inst28_p35),
    .p36(inst28_p36),
    .p37(inst28_p37),
    .p5(inst28_p5),
    .p6(inst28_p6),
    .p7(inst28_p7),
    .p8(inst28_p8),
    .p9(inst28_p9),
    .reset(inst28_reset)
);
comp57 inst29 (
    .clk(inst29_clk),
    .p10(inst29_p10),
    .p11(inst29_p11),
    .p12(inst29_p12),
    .p13(inst29_p13),
    .p14(inst29_p14),
    .p15(inst29_p15),
    .p16(inst29_p16),
    .p17(inst29_p17),
    .p18(inst29_p18),
    .p19(inst29_p19),
    .p20(inst29_p20),
    .p21(inst29_p21),
    .p22(inst29_p22),
    .p23(inst29_p23),
    .p24(inst29_p24),
    .p25(inst29_p25),
    .p26(inst29_p26),
    .p27(inst29_p27),
    .p28(inst29_p28),
    .p29(inst29_p29),
    .p30(inst29_p30),
    .p31(inst29_p31),
    .p32(inst29_p32),
    .p33(inst29_p33),
    .p34(inst29_p34),
    .p35(inst29_p35),
    .p36(inst29_p36),
    .p4(inst29_p4),
    .p5(inst29_p5),
    .p6(inst29_p6),
    .p7(inst29_p7),
    .p8(inst29_p8),
    .p9(inst29_p9),
    .reset(inst29_reset)
);
comp91 inst30 (
    .clk(inst30_clk),
    .p10(inst30_p10),
    .p11(inst30_p11),
    .p12(inst30_p12),
    .p13(inst30_p13),
    .p14(inst30_p14),
    .p15(inst30_p15),
    .p16(inst30_p16),
    .p17(inst30_p17),
    .p18(inst30_p18),
    .p19(inst30_p19),
    .p20(inst30_p20),
    .p21(inst30_p21),
    .p22(inst30_p22),
    .p23(inst30_p23),
    .p24(inst30_p24),
    .p25(inst30_p25),
    .p26(inst30_p26),
    .p27(inst30_p27),
    .p28(inst30_p28),
    .p29(inst30_p29),
    .p30(inst30_p30),
    .p31(inst30_p31),
    .p32(inst30_p32),
    .p33(inst30_p33),
    .p34(inst30_p34),
    .p35(inst30_p35),
    .p36(inst30_p36),
    .p37(inst30_p37),
    .p5(inst30_p5),
    .p6(inst30_p6),
    .p7(inst30_p7),
    .p8(inst30_p8),
    .p9(inst30_p9),
    .reset(inst30_reset)
);
comp57 inst31 (
    .clk(inst31_clk),
    .p10(inst31_p10),
    .p11(inst31_p11),
    .p12(inst31_p12),
    .p13(inst31_p13),
    .p14(inst31_p14),
    .p15(inst31_p15),
    .p16(inst31_p16),
    .p17(inst31_p17),
    .p18(inst31_p18),
    .p19(inst31_p19),
    .p20(inst31_p20),
    .p21(inst31_p21),
    .p22(inst31_p22),
    .p23(inst31_p23),
    .p24(inst31_p24),
    .p25(inst31_p25),
    .p26(inst31_p26),
    .p27(inst31_p27),
    .p28(inst31_p28),
    .p29(inst31_p29),
    .p30(inst31_p30),
    .p31(inst31_p31),
    .p32(inst31_p32),
    .p33(inst31_p33),
    .p34(inst31_p34),
    .p35(inst31_p35),
    .p36(inst31_p36),
    .p4(inst31_p4),
    .p5(inst31_p5),
    .p6(inst31_p6),
    .p7(inst31_p7),
    .p8(inst31_p8),
    .p9(inst31_p9),
    .reset(inst31_reset)
);
comp91 inst32 (
    .clk(inst32_clk),
    .p10(inst32_p10),
    .p11(inst32_p11),
    .p12(inst32_p12),
    .p13(inst32_p13),
    .p14(inst32_p14),
    .p15(inst32_p15),
    .p16(inst32_p16),
    .p17(inst32_p17),
    .p18(inst32_p18),
    .p19(inst32_p19),
    .p20(inst32_p20),
    .p21(inst32_p21),
    .p22(inst32_p22),
    .p23(inst32_p23),
    .p24(inst32_p24),
    .p25(inst32_p25),
    .p26(inst32_p26),
    .p27(inst32_p27),
    .p28(inst32_p28),
    .p29(inst32_p29),
    .p30(inst32_p30),
    .p31(inst32_p31),
    .p32(inst32_p32),
    .p33(inst32_p33),
    .p34(inst32_p34),
    .p35(inst32_p35),
    .p36(inst32_p36),
    .p37(inst32_p37),
    .p5(inst32_p5),
    .p6(inst32_p6),
    .p7(inst32_p7),
    .p8(inst32_p8),
    .p9(inst32_p9),
    .reset(inst32_reset)
);
comp57 inst33 (
    .clk(inst33_clk),
    .p10(inst33_p10),
    .p11(inst33_p11),
    .p12(inst33_p12),
    .p13(inst33_p13),
    .p14(inst33_p14),
    .p15(inst33_p15),
    .p16(inst33_p16),
    .p17(inst33_p17),
    .p18(inst33_p18),
    .p19(inst33_p19),
    .p20(inst33_p20),
    .p21(inst33_p21),
    .p22(inst33_p22),
    .p23(inst33_p23),
    .p24(inst33_p24),
    .p25(inst33_p25),
    .p26(inst33_p26),
    .p27(inst33_p27),
    .p28(inst33_p28),
    .p29(inst33_p29),
    .p30(inst33_p30),
    .p31(inst33_p31),
    .p32(inst33_p32),
    .p33(inst33_p33),
    .p34(inst33_p34),
    .p35(inst33_p35),
    .p36(inst33_p36),
    .p4(inst33_p4),
    .p5(inst33_p5),
    .p6(inst33_p6),
    .p7(inst33_p7),
    .p8(inst33_p8),
    .p9(inst33_p9),
    .reset(inst33_reset)
);
wire _guard0 = 1;
wire _guard1 = ev00__1_0;
wire _guard2 = ev00__1state >= 7'd1;
wire _guard3 = ev00__1state <= 7'd0;
wire _guard4 = _guard2 & _guard3;
wire _guard5 = _guard1 | _guard4;
wire _guard6 = ev00__1_0;
wire _guard7 = ev00__1state >= 7'd1;
wire _guard8 = ev00__1state <= 7'd0;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = _guard6 | _guard9;
wire _guard11 = ev00__1_0;
wire _guard12 = ev00__1state >= 7'd1;
wire _guard13 = ev00__1state <= 7'd0;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = _guard11 | _guard14;
wire _guard16 = ev00__1_0;
wire _guard17 = ev00__1state >= 7'd1;
wire _guard18 = ev00__1state <= 7'd0;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = _guard16 | _guard19;
wire _guard21 = ev00__1_0;
wire _guard22 = ev00__1state >= 7'd1;
wire _guard23 = ev00__1state <= 7'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard21 | _guard24;
wire _guard26 = ev00__1_0;
wire _guard27 = ev00__1state >= 7'd1;
wire _guard28 = ev00__1state <= 7'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard26 | _guard29;
wire _guard31 = ev00__1_0;
wire _guard32 = ev00__1state >= 7'd1;
wire _guard33 = ev00__1state <= 7'd0;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = _guard31 | _guard34;
wire _guard36 = ev00__1_0;
wire _guard37 = ev00__1state >= 7'd1;
wire _guard38 = ev00__1state <= 7'd0;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = _guard36 | _guard39;
wire _guard41 = ev00__1_0;
wire _guard42 = ev00__1state >= 7'd1;
wire _guard43 = ev00__1state <= 7'd0;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = _guard41 | _guard44;
wire _guard46 = ev00__1_0;
wire _guard47 = ev00__1state >= 7'd1;
wire _guard48 = ev00__1state <= 7'd0;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = _guard46 | _guard49;
wire _guard51 = ev00__1_0;
wire _guard52 = ev00__1state >= 7'd1;
wire _guard53 = ev00__1state <= 7'd0;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = _guard51 | _guard54;
wire _guard56 = ev00__1_0;
wire _guard57 = ev00__1state >= 7'd1;
wire _guard58 = ev00__1state <= 7'd0;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = _guard56 | _guard59;
wire _guard61 = ev00__1_0;
wire _guard62 = ev00__1state >= 7'd1;
wire _guard63 = ev00__1state <= 7'd0;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = _guard61 | _guard64;
wire _guard66 = ev00__1_0;
wire _guard67 = ev00__1state >= 7'd1;
wire _guard68 = ev00__1state <= 7'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = _guard66 | _guard69;
wire _guard71 = ev00__1_0;
wire _guard72 = ev00__1state >= 7'd1;
wire _guard73 = ev00__1state <= 7'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard71 | _guard74;
wire _guard76 = ev00__1_0;
wire _guard77 = ev00__1state >= 7'd1;
wire _guard78 = ev00__1state <= 7'd0;
wire _guard79 = _guard77 & _guard78;
wire _guard80 = _guard76 | _guard79;
wire _guard81 = ev00__1_0;
wire _guard82 = ev00__1state >= 7'd1;
wire _guard83 = ev00__1state <= 7'd0;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = _guard81 | _guard84;
wire _guard86 = ev00__1_0;
wire _guard87 = ev00__1state >= 7'd1;
wire _guard88 = ev00__1state <= 7'd0;
wire _guard89 = _guard87 & _guard88;
wire _guard90 = _guard86 | _guard89;
wire _guard91 = ev00__1_0;
wire _guard92 = ev00__1state >= 7'd1;
wire _guard93 = ev00__1state <= 7'd0;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = _guard91 | _guard94;
wire _guard96 = ev00__1_0;
wire _guard97 = ev00__1state >= 7'd1;
wire _guard98 = ev00__1state <= 7'd0;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = _guard96 | _guard99;
wire _guard101 = ev00__1_0;
wire _guard102 = ev00__1state >= 7'd1;
wire _guard103 = ev00__1state <= 7'd0;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = _guard101 | _guard104;
wire _guard106 = ev00__1_0;
wire _guard107 = ev00__1state >= 7'd1;
wire _guard108 = ev00__1state <= 7'd0;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = _guard106 | _guard109;
wire _guard111 = ev00__1_0;
wire _guard112 = ev00__1state >= 7'd1;
wire _guard113 = ev00__1state <= 7'd0;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = _guard111 | _guard114;
wire _guard116 = ev00__1_0;
wire _guard117 = ev00__1state >= 7'd1;
wire _guard118 = ev00__1state <= 7'd0;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = _guard116 | _guard119;
wire _guard121 = ev00__1_0;
wire _guard122 = ev00__1state >= 7'd1;
wire _guard123 = ev00__1state <= 7'd0;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = _guard121 | _guard124;
wire _guard126 = ev00__1_0;
wire _guard127 = ev00__1state >= 7'd1;
wire _guard128 = ev00__1state <= 7'd0;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = _guard126 | _guard129;
wire _guard131 = ev00__1_0;
wire _guard132 = ev00__1state >= 7'd1;
wire _guard133 = ev00__1state <= 7'd0;
wire _guard134 = _guard132 & _guard133;
wire _guard135 = _guard131 | _guard134;
wire _guard136 = ev00__1_0;
wire _guard137 = ev00__1state >= 7'd1;
wire _guard138 = ev00__1state <= 7'd0;
wire _guard139 = _guard137 & _guard138;
wire _guard140 = _guard136 | _guard139;
wire _guard141 = ev00__1_0;
wire _guard142 = ev00__1state >= 7'd1;
wire _guard143 = ev00__1state <= 7'd0;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = _guard141 | _guard144;
wire _guard146 = ev00__1_0;
wire _guard147 = ev00__1state >= 7'd1;
wire _guard148 = ev00__1state <= 7'd0;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = _guard146 | _guard149;
wire _guard151 = ev00__1_0;
wire _guard152 = ev00__1state >= 7'd1;
wire _guard153 = ev00__1state <= 7'd0;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = _guard151 | _guard154;
wire _guard156 = ev00__1_0;
wire _guard157 = ev00__1state >= 7'd1;
wire _guard158 = ev00__1state <= 7'd0;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = _guard156 | _guard159;
wire _guard161 = ev00__0_0;
wire _guard162 = ev00__0state >= 7'd1;
wire _guard163 = ev00__0state <= 7'd127;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = _guard161 | _guard164;
wire _guard166 = ev00__0_0;
wire _guard167 = ev00__0state >= 7'd1;
wire _guard168 = ev00__0state <= 7'd127;
wire _guard169 = _guard167 & _guard168;
wire _guard170 = _guard166 | _guard169;
wire _guard171 = ev00__0_0;
wire _guard172 = ev00__0state >= 7'd1;
wire _guard173 = ev00__0state <= 7'd127;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = _guard171 | _guard174;
wire _guard176 = ev00__0_0;
wire _guard177 = ev00__0state >= 7'd1;
wire _guard178 = ev00__0state <= 7'd127;
wire _guard179 = _guard177 & _guard178;
wire _guard180 = _guard176 | _guard179;
wire _guard181 = ev00__0_0;
wire _guard182 = ev00__0state >= 7'd1;
wire _guard183 = ev00__0state <= 7'd127;
wire _guard184 = _guard182 & _guard183;
wire _guard185 = _guard181 | _guard184;
wire _guard186 = ev00__0_0;
wire _guard187 = ev00__0state >= 7'd1;
wire _guard188 = ev00__0state <= 7'd127;
wire _guard189 = _guard187 & _guard188;
wire _guard190 = _guard186 | _guard189;
wire _guard191 = ev00__0_0;
wire _guard192 = ev00__0state >= 7'd1;
wire _guard193 = ev00__0state <= 7'd127;
wire _guard194 = _guard192 & _guard193;
wire _guard195 = _guard191 | _guard194;
wire _guard196 = ev00__0_0;
wire _guard197 = ev00__0state >= 7'd1;
wire _guard198 = ev00__0state <= 7'd127;
wire _guard199 = _guard197 & _guard198;
wire _guard200 = _guard196 | _guard199;
wire _guard201 = ev00__0_0;
wire _guard202 = ev00__0state >= 7'd1;
wire _guard203 = ev00__0state <= 7'd127;
wire _guard204 = _guard202 & _guard203;
wire _guard205 = _guard201 | _guard204;
wire _guard206 = ev00__0_0;
wire _guard207 = ev00__0state >= 7'd1;
wire _guard208 = ev00__0state <= 7'd127;
wire _guard209 = _guard207 & _guard208;
wire _guard210 = _guard206 | _guard209;
wire _guard211 = ev00__0_0;
wire _guard212 = ev00__0state >= 7'd1;
wire _guard213 = ev00__0state <= 7'd127;
wire _guard214 = _guard212 & _guard213;
wire _guard215 = _guard211 | _guard214;
wire _guard216 = ev00__0_0;
wire _guard217 = ev00__0state >= 7'd1;
wire _guard218 = ev00__0state <= 7'd127;
wire _guard219 = _guard217 & _guard218;
wire _guard220 = _guard216 | _guard219;
wire _guard221 = ev00__0_0;
wire _guard222 = ev00__0state >= 7'd1;
wire _guard223 = ev00__0state <= 7'd127;
wire _guard224 = _guard222 & _guard223;
wire _guard225 = _guard221 | _guard224;
wire _guard226 = ev00__0_0;
wire _guard227 = ev00__0state >= 7'd1;
wire _guard228 = ev00__0state <= 7'd127;
wire _guard229 = _guard227 & _guard228;
wire _guard230 = _guard226 | _guard229;
wire _guard231 = ev00__0_0;
wire _guard232 = ev00__0state >= 7'd1;
wire _guard233 = ev00__0state <= 7'd127;
wire _guard234 = _guard232 & _guard233;
wire _guard235 = _guard231 | _guard234;
wire _guard236 = ev00__0_0;
wire _guard237 = ev00__0state >= 7'd1;
wire _guard238 = ev00__0state <= 7'd127;
wire _guard239 = _guard237 & _guard238;
wire _guard240 = _guard236 | _guard239;
wire _guard241 = ev00__0state >= 7'd95;
wire _guard242 = ev00__0state <= 7'd95;
wire _guard243 = _guard241 & _guard242;
wire _guard244 = ev00__0state >= 7'd32;
wire _guard245 = ev00__0state <= 7'd32;
wire _guard246 = _guard244 & _guard245;
wire _guard247 = ev00__0state >= 7'd32;
wire _guard248 = ev00__0state <= 7'd32;
wire _guard249 = _guard247 & _guard248;
wire _guard250 = ev00__0state >= 7'd32;
wire _guard251 = ev00__0state <= 7'd32;
wire _guard252 = _guard250 & _guard251;
wire _guard253 = ev00__0state >= 7'd32;
wire _guard254 = ev00__0state <= 7'd32;
wire _guard255 = _guard253 & _guard254;
wire _guard256 = ev00__0state >= 7'd32;
wire _guard257 = ev00__0state <= 7'd32;
wire _guard258 = _guard256 & _guard257;
wire _guard259 = ev00__0state >= 7'd32;
wire _guard260 = ev00__0state <= 7'd32;
wire _guard261 = _guard259 & _guard260;
wire _guard262 = ev00__0state >= 7'd32;
wire _guard263 = ev00__0state <= 7'd32;
wire _guard264 = _guard262 & _guard263;
wire _guard265 = ev00__0state >= 7'd32;
wire _guard266 = ev00__0state <= 7'd32;
wire _guard267 = _guard265 & _guard266;
wire _guard268 = ev00__0state >= 7'd32;
wire _guard269 = ev00__0state <= 7'd32;
wire _guard270 = _guard268 & _guard269;
wire _guard271 = ev00__0state >= 7'd32;
wire _guard272 = ev00__0state <= 7'd32;
wire _guard273 = _guard271 & _guard272;
wire _guard274 = ev00__0state >= 7'd32;
wire _guard275 = ev00__0state <= 7'd32;
wire _guard276 = _guard274 & _guard275;
wire _guard277 = ev00__0state >= 7'd32;
wire _guard278 = ev00__0state <= 7'd32;
wire _guard279 = _guard277 & _guard278;
wire _guard280 = ev00__0state >= 7'd32;
wire _guard281 = ev00__0state <= 7'd32;
wire _guard282 = _guard280 & _guard281;
wire _guard283 = ev00__0state >= 7'd32;
wire _guard284 = ev00__0state <= 7'd32;
wire _guard285 = _guard283 & _guard284;
wire _guard286 = ev00__0state >= 7'd32;
wire _guard287 = ev00__0state <= 7'd32;
wire _guard288 = _guard286 & _guard287;
wire _guard289 = ev00__0state >= 7'd32;
wire _guard290 = ev00__0state <= 7'd32;
wire _guard291 = _guard289 & _guard290;
wire _guard292 = ev00__0state >= 7'd32;
wire _guard293 = ev00__0state <= 7'd32;
wire _guard294 = _guard292 & _guard293;
wire _guard295 = ev00__0state >= 7'd32;
wire _guard296 = ev00__0state <= 7'd32;
wire _guard297 = _guard295 & _guard296;
wire _guard298 = ev00__0state >= 7'd32;
wire _guard299 = ev00__0state <= 7'd32;
wire _guard300 = _guard298 & _guard299;
wire _guard301 = ev00__0state >= 7'd32;
wire _guard302 = ev00__0state <= 7'd32;
wire _guard303 = _guard301 & _guard302;
wire _guard304 = ev00__0state >= 7'd32;
wire _guard305 = ev00__0state <= 7'd32;
wire _guard306 = _guard304 & _guard305;
wire _guard307 = ev00__0state >= 7'd32;
wire _guard308 = ev00__0state <= 7'd32;
wire _guard309 = _guard307 & _guard308;
wire _guard310 = ev00__0state >= 7'd32;
wire _guard311 = ev00__0state <= 7'd32;
wire _guard312 = _guard310 & _guard311;
wire _guard313 = ev00__0state >= 7'd32;
wire _guard314 = ev00__0state <= 7'd32;
wire _guard315 = _guard313 & _guard314;
wire _guard316 = ev00__0state >= 7'd32;
wire _guard317 = ev00__0state <= 7'd32;
wire _guard318 = _guard316 & _guard317;
wire _guard319 = ev00__0state >= 7'd32;
wire _guard320 = ev00__0state <= 7'd32;
wire _guard321 = _guard319 & _guard320;
wire _guard322 = ev00__0state >= 7'd32;
wire _guard323 = ev00__0state <= 7'd32;
wire _guard324 = _guard322 & _guard323;
wire _guard325 = ev00__0state >= 7'd32;
wire _guard326 = ev00__0state <= 7'd32;
wire _guard327 = _guard325 & _guard326;
wire _guard328 = ev00__0state >= 7'd32;
wire _guard329 = ev00__0state <= 7'd32;
wire _guard330 = _guard328 & _guard329;
wire _guard331 = ev00__0state >= 7'd32;
wire _guard332 = ev00__0state <= 7'd32;
wire _guard333 = _guard331 & _guard332;
wire _guard334 = ev00__0state >= 7'd32;
wire _guard335 = ev00__0state <= 7'd32;
wire _guard336 = _guard334 & _guard335;
wire _guard337 = ev00__0state >= 7'd32;
wire _guard338 = ev00__0state <= 7'd32;
wire _guard339 = _guard337 & _guard338;
wire _guard340 = ev00__0state >= 7'd62;
wire _guard341 = ev00__0state <= 7'd62;
wire _guard342 = _guard340 & _guard341;
wire _guard343 = ev00__0state >= 7'd62;
wire _guard344 = ev00__0state <= 7'd62;
wire _guard345 = _guard343 & _guard344;
wire _guard346 = ev00__0state >= 7'd62;
wire _guard347 = ev00__0state <= 7'd62;
wire _guard348 = _guard346 & _guard347;
wire _guard349 = ev00__0state >= 7'd62;
wire _guard350 = ev00__0state <= 7'd62;
wire _guard351 = _guard349 & _guard350;
wire _guard352 = ev00__0state >= 7'd62;
wire _guard353 = ev00__0state <= 7'd62;
wire _guard354 = _guard352 & _guard353;
wire _guard355 = ev00__0state >= 7'd62;
wire _guard356 = ev00__0state <= 7'd62;
wire _guard357 = _guard355 & _guard356;
wire _guard358 = ev00__0state >= 7'd62;
wire _guard359 = ev00__0state <= 7'd62;
wire _guard360 = _guard358 & _guard359;
wire _guard361 = ev00__0state >= 7'd62;
wire _guard362 = ev00__0state <= 7'd62;
wire _guard363 = _guard361 & _guard362;
wire _guard364 = ev00__0state >= 7'd62;
wire _guard365 = ev00__0state <= 7'd62;
wire _guard366 = _guard364 & _guard365;
wire _guard367 = ev00__0state >= 7'd62;
wire _guard368 = ev00__0state <= 7'd62;
wire _guard369 = _guard367 & _guard368;
wire _guard370 = ev00__0state >= 7'd62;
wire _guard371 = ev00__0state <= 7'd62;
wire _guard372 = _guard370 & _guard371;
wire _guard373 = ev00__0state >= 7'd62;
wire _guard374 = ev00__0state <= 7'd62;
wire _guard375 = _guard373 & _guard374;
wire _guard376 = ev00__0state >= 7'd62;
wire _guard377 = ev00__0state <= 7'd62;
wire _guard378 = _guard376 & _guard377;
wire _guard379 = ev00__0state >= 7'd62;
wire _guard380 = ev00__0state <= 7'd62;
wire _guard381 = _guard379 & _guard380;
wire _guard382 = ev00__0state >= 7'd62;
wire _guard383 = ev00__0state <= 7'd62;
wire _guard384 = _guard382 & _guard383;
wire _guard385 = ev00__0state >= 7'd62;
wire _guard386 = ev00__0state <= 7'd62;
wire _guard387 = _guard385 & _guard386;
wire _guard388 = ev00__0state >= 7'd62;
wire _guard389 = ev00__0state <= 7'd62;
wire _guard390 = _guard388 & _guard389;
wire _guard391 = ev00__0state >= 7'd62;
wire _guard392 = ev00__0state <= 7'd62;
wire _guard393 = _guard391 & _guard392;
wire _guard394 = ev00__0state >= 7'd62;
wire _guard395 = ev00__0state <= 7'd62;
wire _guard396 = _guard394 & _guard395;
wire _guard397 = ev00__0state >= 7'd62;
wire _guard398 = ev00__0state <= 7'd62;
wire _guard399 = _guard397 & _guard398;
wire _guard400 = ev00__0state >= 7'd62;
wire _guard401 = ev00__0state <= 7'd62;
wire _guard402 = _guard400 & _guard401;
wire _guard403 = ev00__0state >= 7'd62;
wire _guard404 = ev00__0state <= 7'd62;
wire _guard405 = _guard403 & _guard404;
wire _guard406 = ev00__0state >= 7'd62;
wire _guard407 = ev00__0state <= 7'd62;
wire _guard408 = _guard406 & _guard407;
wire _guard409 = ev00__0state >= 7'd62;
wire _guard410 = ev00__0state <= 7'd62;
wire _guard411 = _guard409 & _guard410;
wire _guard412 = ev00__0state >= 7'd62;
wire _guard413 = ev00__0state <= 7'd62;
wire _guard414 = _guard412 & _guard413;
wire _guard415 = ev00__0state >= 7'd62;
wire _guard416 = ev00__0state <= 7'd62;
wire _guard417 = _guard415 & _guard416;
wire _guard418 = ev00__0state >= 7'd62;
wire _guard419 = ev00__0state <= 7'd62;
wire _guard420 = _guard418 & _guard419;
wire _guard421 = ev00__0state >= 7'd62;
wire _guard422 = ev00__0state <= 7'd62;
wire _guard423 = _guard421 & _guard422;
wire _guard424 = ev00__0state >= 7'd62;
wire _guard425 = ev00__0state <= 7'd62;
wire _guard426 = _guard424 & _guard425;
wire _guard427 = ev00__0state >= 7'd62;
wire _guard428 = ev00__0state <= 7'd62;
wire _guard429 = _guard427 & _guard428;
wire _guard430 = ev00__0state >= 7'd62;
wire _guard431 = ev00__0state <= 7'd62;
wire _guard432 = _guard430 & _guard431;
wire _guard433 = ev00__0state >= 7'd62;
wire _guard434 = ev00__0state <= 7'd62;
wire _guard435 = _guard433 & _guard434;
wire _guard436 = ev00__0_0;
wire _guard437 = ev00__0state >= 7'd1;
wire _guard438 = ev00__0state <= 7'd127;
wire _guard439 = _guard437 & _guard438;
wire _guard440 = _guard436 | _guard439;
wire _guard441 = ev00__0_0;
wire _guard442 = ev00__0state >= 7'd1;
wire _guard443 = ev00__0state <= 7'd127;
wire _guard444 = _guard442 & _guard443;
wire _guard445 = _guard441 | _guard444;
wire _guard446 = ev00__0_0;
wire _guard447 = ev00__0state >= 7'd1;
wire _guard448 = ev00__0state <= 7'd127;
wire _guard449 = _guard447 & _guard448;
wire _guard450 = _guard446 | _guard449;
wire _guard451 = ev00__0_0;
wire _guard452 = ev00__0state >= 7'd1;
wire _guard453 = ev00__0state <= 7'd127;
wire _guard454 = _guard452 & _guard453;
wire _guard455 = _guard451 | _guard454;
wire _guard456 = ev00__0_0;
wire _guard457 = ev00__0state >= 7'd1;
wire _guard458 = ev00__0state <= 7'd127;
wire _guard459 = _guard457 & _guard458;
wire _guard460 = _guard456 | _guard459;
wire _guard461 = ev00__0_0;
wire _guard462 = ev00__0state >= 7'd1;
wire _guard463 = ev00__0state <= 7'd127;
wire _guard464 = _guard462 & _guard463;
wire _guard465 = _guard461 | _guard464;
wire _guard466 = ev00__0_0;
wire _guard467 = ev00__0state >= 7'd1;
wire _guard468 = ev00__0state <= 7'd127;
wire _guard469 = _guard467 & _guard468;
wire _guard470 = _guard466 | _guard469;
wire _guard471 = ev00__0_0;
wire _guard472 = ev00__0state >= 7'd1;
wire _guard473 = ev00__0state <= 7'd127;
wire _guard474 = _guard472 & _guard473;
wire _guard475 = _guard471 | _guard474;
wire _guard476 = ev00__0_0;
wire _guard477 = ev00__0state >= 7'd1;
wire _guard478 = ev00__0state <= 7'd127;
wire _guard479 = _guard477 & _guard478;
wire _guard480 = _guard476 | _guard479;
wire _guard481 = ev00__0_0;
wire _guard482 = ev00__0state >= 7'd1;
wire _guard483 = ev00__0state <= 7'd127;
wire _guard484 = _guard482 & _guard483;
wire _guard485 = _guard481 | _guard484;
wire _guard486 = ev00__0_0;
wire _guard487 = ev00__0state >= 7'd1;
wire _guard488 = ev00__0state <= 7'd127;
wire _guard489 = _guard487 & _guard488;
wire _guard490 = _guard486 | _guard489;
wire _guard491 = ev00__0_0;
wire _guard492 = ev00__0state >= 7'd1;
wire _guard493 = ev00__0state <= 7'd127;
wire _guard494 = _guard492 & _guard493;
wire _guard495 = _guard491 | _guard494;
wire _guard496 = ev00__0_0;
wire _guard497 = ev00__0state >= 7'd1;
wire _guard498 = ev00__0state <= 7'd127;
wire _guard499 = _guard497 & _guard498;
wire _guard500 = _guard496 | _guard499;
wire _guard501 = ev00__0_0;
wire _guard502 = ev00__0state >= 7'd1;
wire _guard503 = ev00__0state <= 7'd127;
wire _guard504 = _guard502 & _guard503;
wire _guard505 = _guard501 | _guard504;
wire _guard506 = ev00__0_0;
wire _guard507 = ev00__0state >= 7'd1;
wire _guard508 = ev00__0state <= 7'd127;
wire _guard509 = _guard507 & _guard508;
wire _guard510 = _guard506 | _guard509;
wire _guard511 = ev00__0_0;
wire _guard512 = ev00__0state >= 7'd1;
wire _guard513 = ev00__0state <= 7'd127;
wire _guard514 = _guard512 & _guard513;
wire _guard515 = _guard511 | _guard514;
wire _guard516 = ev00__0state >= 7'd30;
wire _guard517 = ev00__0state <= 7'd30;
wire _guard518 = _guard516 & _guard517;
wire _guard519 = ev00__0state >= 7'd30;
wire _guard520 = ev00__0state <= 7'd30;
wire _guard521 = _guard519 & _guard520;
wire _guard522 = ev00__0state >= 7'd30;
wire _guard523 = ev00__0state <= 7'd30;
wire _guard524 = _guard522 & _guard523;
wire _guard525 = ev00__0state >= 7'd30;
wire _guard526 = ev00__0state <= 7'd30;
wire _guard527 = _guard525 & _guard526;
wire _guard528 = ev00__0state >= 7'd30;
wire _guard529 = ev00__0state <= 7'd30;
wire _guard530 = _guard528 & _guard529;
wire _guard531 = ev00__0state >= 7'd30;
wire _guard532 = ev00__0state <= 7'd30;
wire _guard533 = _guard531 & _guard532;
wire _guard534 = ev00__0state >= 7'd30;
wire _guard535 = ev00__0state <= 7'd30;
wire _guard536 = _guard534 & _guard535;
wire _guard537 = ev00__0state >= 7'd30;
wire _guard538 = ev00__0state <= 7'd30;
wire _guard539 = _guard537 & _guard538;
wire _guard540 = ev00__0state >= 7'd30;
wire _guard541 = ev00__0state <= 7'd30;
wire _guard542 = _guard540 & _guard541;
wire _guard543 = ev00__0state >= 7'd30;
wire _guard544 = ev00__0state <= 7'd30;
wire _guard545 = _guard543 & _guard544;
wire _guard546 = ev00__0state >= 7'd30;
wire _guard547 = ev00__0state <= 7'd30;
wire _guard548 = _guard546 & _guard547;
wire _guard549 = ev00__0state >= 7'd30;
wire _guard550 = ev00__0state <= 7'd30;
wire _guard551 = _guard549 & _guard550;
wire _guard552 = ev00__0state >= 7'd30;
wire _guard553 = ev00__0state <= 7'd30;
wire _guard554 = _guard552 & _guard553;
wire _guard555 = ev00__0state >= 7'd30;
wire _guard556 = ev00__0state <= 7'd30;
wire _guard557 = _guard555 & _guard556;
wire _guard558 = ev00__0state >= 7'd30;
wire _guard559 = ev00__0state <= 7'd30;
wire _guard560 = _guard558 & _guard559;
wire _guard561 = ev00__0state >= 7'd30;
wire _guard562 = ev00__0state <= 7'd30;
wire _guard563 = _guard561 & _guard562;
wire _guard564 = ev00__0state >= 7'd30;
wire _guard565 = ev00__0state <= 7'd30;
wire _guard566 = _guard564 & _guard565;
wire _guard567 = ev00__0state >= 7'd30;
wire _guard568 = ev00__0state <= 7'd30;
wire _guard569 = _guard567 & _guard568;
wire _guard570 = ev00__0state >= 7'd30;
wire _guard571 = ev00__0state <= 7'd30;
wire _guard572 = _guard570 & _guard571;
wire _guard573 = ev00__0state >= 7'd30;
wire _guard574 = ev00__0state <= 7'd30;
wire _guard575 = _guard573 & _guard574;
wire _guard576 = ev00__0state >= 7'd30;
wire _guard577 = ev00__0state <= 7'd30;
wire _guard578 = _guard576 & _guard577;
wire _guard579 = ev00__0state >= 7'd30;
wire _guard580 = ev00__0state <= 7'd30;
wire _guard581 = _guard579 & _guard580;
wire _guard582 = ev00__0state >= 7'd30;
wire _guard583 = ev00__0state <= 7'd30;
wire _guard584 = _guard582 & _guard583;
wire _guard585 = ev00__0state >= 7'd30;
wire _guard586 = ev00__0state <= 7'd30;
wire _guard587 = _guard585 & _guard586;
wire _guard588 = ev00__0state >= 7'd30;
wire _guard589 = ev00__0state <= 7'd30;
wire _guard590 = _guard588 & _guard589;
wire _guard591 = ev00__0state >= 7'd30;
wire _guard592 = ev00__0state <= 7'd30;
wire _guard593 = _guard591 & _guard592;
wire _guard594 = ev00__0state >= 7'd30;
wire _guard595 = ev00__0state <= 7'd30;
wire _guard596 = _guard594 & _guard595;
wire _guard597 = ev00__0state >= 7'd30;
wire _guard598 = ev00__0state <= 7'd30;
wire _guard599 = _guard597 & _guard598;
wire _guard600 = ev00__0state >= 7'd30;
wire _guard601 = ev00__0state <= 7'd30;
wire _guard602 = _guard600 & _guard601;
wire _guard603 = ev00__0state >= 7'd30;
wire _guard604 = ev00__0state <= 7'd30;
wire _guard605 = _guard603 & _guard604;
wire _guard606 = ev00__0state >= 7'd30;
wire _guard607 = ev00__0state <= 7'd30;
wire _guard608 = _guard606 & _guard607;
wire _guard609 = ev00__0state >= 7'd30;
wire _guard610 = ev00__0state <= 7'd30;
wire _guard611 = _guard609 & _guard610;
wire _guard612 = ev00__0state >= 7'd96;
wire _guard613 = ev00__0state <= 7'd96;
wire _guard614 = _guard612 & _guard613;
wire _guard615 = ev00__0state >= 7'd127;
wire _guard616 = ev00__0state <= 7'd127;
wire _guard617 = _guard615 & _guard616;
wire _guard618 = ev00__0state >= 7'd127;
wire _guard619 = ev00__0state <= 7'd127;
wire _guard620 = _guard618 & _guard619;
wire _guard621 = ev00__0state >= 7'd127;
wire _guard622 = ev00__0state <= 7'd127;
wire _guard623 = _guard621 & _guard622;
wire _guard624 = ev00__0state >= 7'd127;
wire _guard625 = ev00__0state <= 7'd127;
wire _guard626 = _guard624 & _guard625;
wire _guard627 = ev00__0state >= 7'd127;
wire _guard628 = ev00__0state <= 7'd127;
wire _guard629 = _guard627 & _guard628;
wire _guard630 = ev00__0state >= 7'd127;
wire _guard631 = ev00__0state <= 7'd127;
wire _guard632 = _guard630 & _guard631;
wire _guard633 = ev00__0state >= 7'd127;
wire _guard634 = ev00__0state <= 7'd127;
wire _guard635 = _guard633 & _guard634;
wire _guard636 = ev00__0state >= 7'd127;
wire _guard637 = ev00__0state <= 7'd127;
wire _guard638 = _guard636 & _guard637;
wire _guard639 = ev00__0state >= 7'd127;
wire _guard640 = ev00__0state <= 7'd127;
wire _guard641 = _guard639 & _guard640;
wire _guard642 = ev00__0state >= 7'd127;
wire _guard643 = ev00__0state <= 7'd127;
wire _guard644 = _guard642 & _guard643;
wire _guard645 = ev00__0state >= 7'd127;
wire _guard646 = ev00__0state <= 7'd127;
wire _guard647 = _guard645 & _guard646;
wire _guard648 = ev00__0state >= 7'd127;
wire _guard649 = ev00__0state <= 7'd127;
wire _guard650 = _guard648 & _guard649;
wire _guard651 = ev00__0state >= 7'd127;
wire _guard652 = ev00__0state <= 7'd127;
wire _guard653 = _guard651 & _guard652;
wire _guard654 = ev00__0state >= 7'd127;
wire _guard655 = ev00__0state <= 7'd127;
wire _guard656 = _guard654 & _guard655;
wire _guard657 = ev00__0state >= 7'd127;
wire _guard658 = ev00__0state <= 7'd127;
wire _guard659 = _guard657 & _guard658;
wire _guard660 = ev00__0state >= 7'd127;
wire _guard661 = ev00__0state <= 7'd127;
wire _guard662 = _guard660 & _guard661;
wire _guard663 = ev00__0state >= 7'd127;
wire _guard664 = ev00__0state <= 7'd127;
wire _guard665 = _guard663 & _guard664;
wire _guard666 = ev00__0state >= 7'd127;
wire _guard667 = ev00__0state <= 7'd127;
wire _guard668 = _guard666 & _guard667;
wire _guard669 = ev00__0state >= 7'd127;
wire _guard670 = ev00__0state <= 7'd127;
wire _guard671 = _guard669 & _guard670;
wire _guard672 = ev00__0state >= 7'd127;
wire _guard673 = ev00__0state <= 7'd127;
wire _guard674 = _guard672 & _guard673;
wire _guard675 = ev00__0state >= 7'd127;
wire _guard676 = ev00__0state <= 7'd127;
wire _guard677 = _guard675 & _guard676;
wire _guard678 = ev00__0state >= 7'd127;
wire _guard679 = ev00__0state <= 7'd127;
wire _guard680 = _guard678 & _guard679;
wire _guard681 = ev00__0state >= 7'd127;
wire _guard682 = ev00__0state <= 7'd127;
wire _guard683 = _guard681 & _guard682;
wire _guard684 = ev00__0state >= 7'd127;
wire _guard685 = ev00__0state <= 7'd127;
wire _guard686 = _guard684 & _guard685;
wire _guard687 = ev00__0state >= 7'd127;
wire _guard688 = ev00__0state <= 7'd127;
wire _guard689 = _guard687 & _guard688;
wire _guard690 = ev00__0state >= 7'd127;
wire _guard691 = ev00__0state <= 7'd127;
wire _guard692 = _guard690 & _guard691;
wire _guard693 = ev00__0state >= 7'd127;
wire _guard694 = ev00__0state <= 7'd127;
wire _guard695 = _guard693 & _guard694;
wire _guard696 = ev00__0state >= 7'd127;
wire _guard697 = ev00__0state <= 7'd127;
wire _guard698 = _guard696 & _guard697;
wire _guard699 = ev00__0state >= 7'd127;
wire _guard700 = ev00__0state <= 7'd127;
wire _guard701 = _guard699 & _guard700;
wire _guard702 = ev00__0state >= 7'd127;
wire _guard703 = ev00__0state <= 7'd127;
wire _guard704 = _guard702 & _guard703;
wire _guard705 = ev00__0state >= 7'd127;
wire _guard706 = ev00__0state <= 7'd127;
wire _guard707 = _guard705 & _guard706;
wire _guard708 = ev00__0state >= 7'd127;
wire _guard709 = ev00__0state <= 7'd127;
wire _guard710 = _guard708 & _guard709;
wire _guard711 = ev00__0_0;
wire _guard712 = ev00__0state >= 7'd1;
wire _guard713 = ev00__0state <= 7'd0;
wire _guard714 = _guard712 & _guard713;
wire _guard715 = _guard711 | _guard714;
wire _guard716 = ev00__0_0;
wire _guard717 = ev00__0state >= 7'd1;
wire _guard718 = ev00__0state <= 7'd0;
wire _guard719 = _guard717 & _guard718;
wire _guard720 = _guard716 | _guard719;
wire _guard721 = ev00__0_0;
wire _guard722 = ev00__0state >= 7'd1;
wire _guard723 = ev00__0state <= 7'd0;
wire _guard724 = _guard722 & _guard723;
wire _guard725 = _guard721 | _guard724;
wire _guard726 = ev00__0_0;
wire _guard727 = ev00__0state >= 7'd1;
wire _guard728 = ev00__0state <= 7'd0;
wire _guard729 = _guard727 & _guard728;
wire _guard730 = _guard726 | _guard729;
wire _guard731 = ev00__0_0;
wire _guard732 = ev00__0state >= 7'd1;
wire _guard733 = ev00__0state <= 7'd0;
wire _guard734 = _guard732 & _guard733;
wire _guard735 = _guard731 | _guard734;
wire _guard736 = ev00__0_0;
wire _guard737 = ev00__0state >= 7'd1;
wire _guard738 = ev00__0state <= 7'd0;
wire _guard739 = _guard737 & _guard738;
wire _guard740 = _guard736 | _guard739;
wire _guard741 = ev00__0_0;
wire _guard742 = ev00__0state >= 7'd1;
wire _guard743 = ev00__0state <= 7'd0;
wire _guard744 = _guard742 & _guard743;
wire _guard745 = _guard741 | _guard744;
wire _guard746 = ev00__0_0;
wire _guard747 = ev00__0state >= 7'd1;
wire _guard748 = ev00__0state <= 7'd0;
wire _guard749 = _guard747 & _guard748;
wire _guard750 = _guard746 | _guard749;
wire _guard751 = ev00__0_0;
wire _guard752 = ev00__0state >= 7'd1;
wire _guard753 = ev00__0state <= 7'd0;
wire _guard754 = _guard752 & _guard753;
wire _guard755 = _guard751 | _guard754;
wire _guard756 = ev00__0_0;
wire _guard757 = ev00__0state >= 7'd1;
wire _guard758 = ev00__0state <= 7'd0;
wire _guard759 = _guard757 & _guard758;
wire _guard760 = _guard756 | _guard759;
wire _guard761 = ev00__0_0;
wire _guard762 = ev00__0state >= 7'd1;
wire _guard763 = ev00__0state <= 7'd0;
wire _guard764 = _guard762 & _guard763;
wire _guard765 = _guard761 | _guard764;
wire _guard766 = ev00__0_0;
wire _guard767 = ev00__0state >= 7'd1;
wire _guard768 = ev00__0state <= 7'd0;
wire _guard769 = _guard767 & _guard768;
wire _guard770 = _guard766 | _guard769;
wire _guard771 = ev00__0_0;
wire _guard772 = ev00__0state >= 7'd1;
wire _guard773 = ev00__0state <= 7'd0;
wire _guard774 = _guard772 & _guard773;
wire _guard775 = _guard771 | _guard774;
wire _guard776 = ev00__0_0;
wire _guard777 = ev00__0state >= 7'd1;
wire _guard778 = ev00__0state <= 7'd0;
wire _guard779 = _guard777 & _guard778;
wire _guard780 = _guard776 | _guard779;
wire _guard781 = ev00__0_0;
wire _guard782 = ev00__0state >= 7'd1;
wire _guard783 = ev00__0state <= 7'd0;
wire _guard784 = _guard782 & _guard783;
wire _guard785 = _guard781 | _guard784;
wire _guard786 = ev00__0_0;
wire _guard787 = ev00__0state >= 7'd1;
wire _guard788 = ev00__0state <= 7'd0;
wire _guard789 = _guard787 & _guard788;
wire _guard790 = _guard786 | _guard789;
wire _guard791 = ev00__0_0;
wire _guard792 = ev00__0state >= 7'd1;
wire _guard793 = ev00__0state <= 7'd0;
wire _guard794 = _guard792 & _guard793;
wire _guard795 = _guard791 | _guard794;
wire _guard796 = ev00__0_0;
wire _guard797 = ev00__0state >= 7'd1;
wire _guard798 = ev00__0state <= 7'd0;
wire _guard799 = _guard797 & _guard798;
wire _guard800 = _guard796 | _guard799;
wire _guard801 = ev00__0_0;
wire _guard802 = ev00__0state >= 7'd1;
wire _guard803 = ev00__0state <= 7'd0;
wire _guard804 = _guard802 & _guard803;
wire _guard805 = _guard801 | _guard804;
wire _guard806 = ev00__0_0;
wire _guard807 = ev00__0state >= 7'd1;
wire _guard808 = ev00__0state <= 7'd0;
wire _guard809 = _guard807 & _guard808;
wire _guard810 = _guard806 | _guard809;
wire _guard811 = ev00__0_0;
wire _guard812 = ev00__0state >= 7'd1;
wire _guard813 = ev00__0state <= 7'd0;
wire _guard814 = _guard812 & _guard813;
wire _guard815 = _guard811 | _guard814;
wire _guard816 = ev00__0_0;
wire _guard817 = ev00__0state >= 7'd1;
wire _guard818 = ev00__0state <= 7'd0;
wire _guard819 = _guard817 & _guard818;
wire _guard820 = _guard816 | _guard819;
wire _guard821 = ev00__0_0;
wire _guard822 = ev00__0state >= 7'd1;
wire _guard823 = ev00__0state <= 7'd0;
wire _guard824 = _guard822 & _guard823;
wire _guard825 = _guard821 | _guard824;
wire _guard826 = ev00__0_0;
wire _guard827 = ev00__0state >= 7'd1;
wire _guard828 = ev00__0state <= 7'd0;
wire _guard829 = _guard827 & _guard828;
wire _guard830 = _guard826 | _guard829;
wire _guard831 = ev00__0_0;
wire _guard832 = ev00__0state >= 7'd1;
wire _guard833 = ev00__0state <= 7'd0;
wire _guard834 = _guard832 & _guard833;
wire _guard835 = _guard831 | _guard834;
wire _guard836 = ev00__0_0;
wire _guard837 = ev00__0state >= 7'd1;
wire _guard838 = ev00__0state <= 7'd0;
wire _guard839 = _guard837 & _guard838;
wire _guard840 = _guard836 | _guard839;
wire _guard841 = ev00__0_0;
wire _guard842 = ev00__0state >= 7'd1;
wire _guard843 = ev00__0state <= 7'd0;
wire _guard844 = _guard842 & _guard843;
wire _guard845 = _guard841 | _guard844;
wire _guard846 = ev00__0_0;
wire _guard847 = ev00__0state >= 7'd1;
wire _guard848 = ev00__0state <= 7'd0;
wire _guard849 = _guard847 & _guard848;
wire _guard850 = _guard846 | _guard849;
wire _guard851 = ev00__0_0;
wire _guard852 = ev00__0state >= 7'd1;
wire _guard853 = ev00__0state <= 7'd0;
wire _guard854 = _guard852 & _guard853;
wire _guard855 = _guard851 | _guard854;
wire _guard856 = ev00__0_0;
wire _guard857 = ev00__0state >= 7'd1;
wire _guard858 = ev00__0state <= 7'd0;
wire _guard859 = _guard857 & _guard858;
wire _guard860 = _guard856 | _guard859;
wire _guard861 = ev00__0_0;
wire _guard862 = ev00__0state >= 7'd1;
wire _guard863 = ev00__0state <= 7'd0;
wire _guard864 = _guard862 & _guard863;
wire _guard865 = _guard861 | _guard864;
wire _guard866 = ev00__0_0;
wire _guard867 = ev00__0state >= 7'd1;
wire _guard868 = ev00__0state <= 7'd0;
wire _guard869 = _guard867 & _guard868;
wire _guard870 = _guard866 | _guard869;
wire _guard871 = ev00__0state >= 7'd127;
wire _guard872 = ev00__0state <= 7'd127;
wire _guard873 = _guard871 & _guard872;
wire _guard874 = ev00__0state >= 7'd64;
wire _guard875 = ev00__0state <= 7'd64;
wire _guard876 = _guard874 & _guard875;
wire _guard877 = ev00__0state >= 7'd63;
wire _guard878 = ev00__0state <= 7'd63;
wire _guard879 = _guard877 & _guard878;
wire _guard880 = ev00__0state >= 7'd63;
wire _guard881 = ev00__0state <= 7'd63;
wire _guard882 = _guard880 & _guard881;
wire _guard883 = ev00__0state >= 7'd63;
wire _guard884 = ev00__0state <= 7'd63;
wire _guard885 = _guard883 & _guard884;
wire _guard886 = ev00__0state >= 7'd63;
wire _guard887 = ev00__0state <= 7'd63;
wire _guard888 = _guard886 & _guard887;
wire _guard889 = ev00__0state >= 7'd63;
wire _guard890 = ev00__0state <= 7'd63;
wire _guard891 = _guard889 & _guard890;
wire _guard892 = ev00__0state >= 7'd63;
wire _guard893 = ev00__0state <= 7'd63;
wire _guard894 = _guard892 & _guard893;
wire _guard895 = ev00__0state >= 7'd63;
wire _guard896 = ev00__0state <= 7'd63;
wire _guard897 = _guard895 & _guard896;
wire _guard898 = ev00__0state >= 7'd63;
wire _guard899 = ev00__0state <= 7'd63;
wire _guard900 = _guard898 & _guard899;
wire _guard901 = ev00__0state >= 7'd63;
wire _guard902 = ev00__0state <= 7'd63;
wire _guard903 = _guard901 & _guard902;
wire _guard904 = ev00__0state >= 7'd63;
wire _guard905 = ev00__0state <= 7'd63;
wire _guard906 = _guard904 & _guard905;
wire _guard907 = ev00__0state >= 7'd63;
wire _guard908 = ev00__0state <= 7'd63;
wire _guard909 = _guard907 & _guard908;
wire _guard910 = ev00__0state >= 7'd63;
wire _guard911 = ev00__0state <= 7'd63;
wire _guard912 = _guard910 & _guard911;
wire _guard913 = ev00__0state >= 7'd63;
wire _guard914 = ev00__0state <= 7'd63;
wire _guard915 = _guard913 & _guard914;
wire _guard916 = ev00__0state >= 7'd63;
wire _guard917 = ev00__0state <= 7'd63;
wire _guard918 = _guard916 & _guard917;
wire _guard919 = ev00__0state >= 7'd63;
wire _guard920 = ev00__0state <= 7'd63;
wire _guard921 = _guard919 & _guard920;
wire _guard922 = ev00__0state >= 7'd63;
wire _guard923 = ev00__0state <= 7'd63;
wire _guard924 = _guard922 & _guard923;
wire _guard925 = ev00__0state >= 7'd63;
wire _guard926 = ev00__0state <= 7'd63;
wire _guard927 = _guard925 & _guard926;
wire _guard928 = ev00__0state >= 7'd63;
wire _guard929 = ev00__0state <= 7'd63;
wire _guard930 = _guard928 & _guard929;
wire _guard931 = ev00__0state >= 7'd63;
wire _guard932 = ev00__0state <= 7'd63;
wire _guard933 = _guard931 & _guard932;
wire _guard934 = ev00__0state >= 7'd63;
wire _guard935 = ev00__0state <= 7'd63;
wire _guard936 = _guard934 & _guard935;
wire _guard937 = ev00__0state >= 7'd63;
wire _guard938 = ev00__0state <= 7'd63;
wire _guard939 = _guard937 & _guard938;
wire _guard940 = ev00__0state >= 7'd63;
wire _guard941 = ev00__0state <= 7'd63;
wire _guard942 = _guard940 & _guard941;
wire _guard943 = ev00__0state >= 7'd63;
wire _guard944 = ev00__0state <= 7'd63;
wire _guard945 = _guard943 & _guard944;
wire _guard946 = ev00__0state >= 7'd63;
wire _guard947 = ev00__0state <= 7'd63;
wire _guard948 = _guard946 & _guard947;
wire _guard949 = ev00__0state >= 7'd63;
wire _guard950 = ev00__0state <= 7'd63;
wire _guard951 = _guard949 & _guard950;
wire _guard952 = ev00__0state >= 7'd63;
wire _guard953 = ev00__0state <= 7'd63;
wire _guard954 = _guard952 & _guard953;
wire _guard955 = ev00__0state >= 7'd63;
wire _guard956 = ev00__0state <= 7'd63;
wire _guard957 = _guard955 & _guard956;
wire _guard958 = ev00__0state >= 7'd63;
wire _guard959 = ev00__0state <= 7'd63;
wire _guard960 = _guard958 & _guard959;
wire _guard961 = ev00__0state >= 7'd63;
wire _guard962 = ev00__0state <= 7'd63;
wire _guard963 = _guard961 & _guard962;
wire _guard964 = ev00__0state >= 7'd63;
wire _guard965 = ev00__0state <= 7'd63;
wire _guard966 = _guard964 & _guard965;
wire _guard967 = ev00__0state >= 7'd63;
wire _guard968 = ev00__0state <= 7'd63;
wire _guard969 = _guard967 & _guard968;
wire _guard970 = ev00__0state >= 7'd63;
wire _guard971 = ev00__0state <= 7'd63;
wire _guard972 = _guard970 & _guard971;
wire _guard973 = ev00__0_0;
wire _guard974 = ev00__0state >= 7'd1;
wire _guard975 = ev00__0state <= 7'd0;
wire _guard976 = _guard974 & _guard975;
wire _guard977 = _guard973 | _guard976;
wire _guard978 = ev00__0state >= 7'd30;
wire _guard979 = ev00__0state <= 7'd30;
wire _guard980 = _guard978 & _guard979;
wire _guard981 = _guard977 | _guard980;
wire _guard982 = ev00__0state >= 7'd32;
wire _guard983 = ev00__0state <= 7'd32;
wire _guard984 = _guard982 & _guard983;
wire _guard985 = _guard981 | _guard984;
wire _guard986 = ev00__0state >= 7'd62;
wire _guard987 = ev00__0state <= 7'd62;
wire _guard988 = _guard986 & _guard987;
wire _guard989 = _guard985 | _guard988;
wire _guard990 = ev00__0state >= 7'd64;
wire _guard991 = ev00__0state <= 7'd64;
wire _guard992 = _guard990 & _guard991;
wire _guard993 = _guard989 | _guard992;
wire _guard994 = ev00__0state >= 7'd94;
wire _guard995 = ev00__0state <= 7'd94;
wire _guard996 = _guard994 & _guard995;
wire _guard997 = _guard993 | _guard996;
wire _guard998 = ev00__0state >= 7'd96;
wire _guard999 = ev00__0state <= 7'd96;
wire _guard1000 = _guard998 & _guard999;
wire _guard1001 = _guard997 | _guard1000;
wire _guard1002 = ev00__0state >= 7'd126;
wire _guard1003 = ev00__0state <= 7'd126;
wire _guard1004 = _guard1002 & _guard1003;
wire _guard1005 = _guard1001 | _guard1004;
wire _guard1006 = ev00__0state >= 7'd32;
wire _guard1007 = ev00__0state <= 7'd32;
wire _guard1008 = _guard1006 & _guard1007;
wire _guard1009 = ev00__0state >= 7'd62;
wire _guard1010 = ev00__0state <= 7'd62;
wire _guard1011 = _guard1009 & _guard1010;
wire _guard1012 = ev00__0state >= 7'd30;
wire _guard1013 = ev00__0state <= 7'd30;
wire _guard1014 = _guard1012 & _guard1013;
wire _guard1015 = ev00__0state >= 7'd126;
wire _guard1016 = ev00__0state <= 7'd126;
wire _guard1017 = _guard1015 & _guard1016;
wire _guard1018 = ev00__0state >= 7'd96;
wire _guard1019 = ev00__0state <= 7'd96;
wire _guard1020 = _guard1018 & _guard1019;
wire _guard1021 = ev00__0state >= 7'd64;
wire _guard1022 = ev00__0state <= 7'd64;
wire _guard1023 = _guard1021 & _guard1022;
wire _guard1024 = ev00__0state >= 7'd94;
wire _guard1025 = ev00__0state <= 7'd94;
wire _guard1026 = _guard1024 & _guard1025;
wire _guard1027 = ev00__0_0;
wire _guard1028 = ev00__0state >= 7'd1;
wire _guard1029 = ev00__0state <= 7'd0;
wire _guard1030 = _guard1028 & _guard1029;
wire _guard1031 = _guard1027 | _guard1030;
wire _guard1032 = ev00__0state >= 7'd63;
wire _guard1033 = ev00__0state <= 7'd63;
wire _guard1034 = _guard1032 & _guard1033;
wire _guard1035 = ev00__0state >= 7'd95;
wire _guard1036 = ev00__0state <= 7'd95;
wire _guard1037 = _guard1035 & _guard1036;
wire _guard1038 = ev00__0state >= 7'd127;
wire _guard1039 = ev00__0state <= 7'd127;
wire _guard1040 = _guard1038 & _guard1039;
wire _guard1041 = ev00__0state >= 7'd63;
wire _guard1042 = ev00__0state <= 7'd63;
wire _guard1043 = _guard1041 & _guard1042;
wire _guard1044 = ev00__0state >= 7'd31;
wire _guard1045 = ev00__0state <= 7'd31;
wire _guard1046 = _guard1044 & _guard1045;
wire _guard1047 = ev00__0state >= 7'd95;
wire _guard1048 = ev00__0state <= 7'd95;
wire _guard1049 = _guard1047 & _guard1048;
wire _guard1050 = ev00__0state >= 7'd127;
wire _guard1051 = ev00__0state <= 7'd127;
wire _guard1052 = _guard1050 & _guard1051;
wire _guard1053 = ev00__0state >= 7'd63;
wire _guard1054 = ev00__0state <= 7'd63;
wire _guard1055 = _guard1053 & _guard1054;
wire _guard1056 = ev00__0state >= 7'd31;
wire _guard1057 = ev00__0state <= 7'd31;
wire _guard1058 = _guard1056 & _guard1057;
wire _guard1059 = ev00__0state >= 7'd95;
wire _guard1060 = ev00__0state <= 7'd95;
wire _guard1061 = _guard1059 & _guard1060;
wire _guard1062 = ev00__0state >= 7'd127;
wire _guard1063 = ev00__0state <= 7'd127;
wire _guard1064 = _guard1062 & _guard1063;
wire _guard1065 = ev00__0state >= 7'd63;
wire _guard1066 = ev00__0state <= 7'd63;
wire _guard1067 = _guard1065 & _guard1066;
wire _guard1068 = ev00__0state >= 7'd31;
wire _guard1069 = ev00__0state <= 7'd31;
wire _guard1070 = _guard1068 & _guard1069;
wire _guard1071 = ev00__0state >= 7'd95;
wire _guard1072 = ev00__0state <= 7'd95;
wire _guard1073 = _guard1071 & _guard1072;
wire _guard1074 = ev00__0state >= 7'd127;
wire _guard1075 = ev00__0state <= 7'd127;
wire _guard1076 = _guard1074 & _guard1075;
wire _guard1077 = ev00__0state >= 7'd63;
wire _guard1078 = ev00__0state <= 7'd63;
wire _guard1079 = _guard1077 & _guard1078;
wire _guard1080 = ev00__0state >= 7'd31;
wire _guard1081 = ev00__0state <= 7'd31;
wire _guard1082 = _guard1080 & _guard1081;
wire _guard1083 = ev00__0state >= 7'd95;
wire _guard1084 = ev00__0state <= 7'd95;
wire _guard1085 = _guard1083 & _guard1084;
wire _guard1086 = ev00__0state >= 7'd127;
wire _guard1087 = ev00__0state <= 7'd127;
wire _guard1088 = _guard1086 & _guard1087;
wire _guard1089 = ev00__0state >= 7'd63;
wire _guard1090 = ev00__0state <= 7'd63;
wire _guard1091 = _guard1089 & _guard1090;
wire _guard1092 = ev00__0state >= 7'd31;
wire _guard1093 = ev00__0state <= 7'd31;
wire _guard1094 = _guard1092 & _guard1093;
wire _guard1095 = ev00__0state >= 7'd95;
wire _guard1096 = ev00__0state <= 7'd95;
wire _guard1097 = _guard1095 & _guard1096;
wire _guard1098 = ev00__0state >= 7'd127;
wire _guard1099 = ev00__0state <= 7'd127;
wire _guard1100 = _guard1098 & _guard1099;
wire _guard1101 = ev00__0state >= 7'd63;
wire _guard1102 = ev00__0state <= 7'd63;
wire _guard1103 = _guard1101 & _guard1102;
wire _guard1104 = ev00__0state >= 7'd31;
wire _guard1105 = ev00__0state <= 7'd31;
wire _guard1106 = _guard1104 & _guard1105;
wire _guard1107 = ev00__0state >= 7'd95;
wire _guard1108 = ev00__0state <= 7'd95;
wire _guard1109 = _guard1107 & _guard1108;
wire _guard1110 = ev00__0state >= 7'd127;
wire _guard1111 = ev00__0state <= 7'd127;
wire _guard1112 = _guard1110 & _guard1111;
wire _guard1113 = ev00__0state >= 7'd63;
wire _guard1114 = ev00__0state <= 7'd63;
wire _guard1115 = _guard1113 & _guard1114;
wire _guard1116 = ev00__0state >= 7'd31;
wire _guard1117 = ev00__0state <= 7'd31;
wire _guard1118 = _guard1116 & _guard1117;
wire _guard1119 = ev00__0state >= 7'd95;
wire _guard1120 = ev00__0state <= 7'd95;
wire _guard1121 = _guard1119 & _guard1120;
wire _guard1122 = ev00__0state >= 7'd127;
wire _guard1123 = ev00__0state <= 7'd127;
wire _guard1124 = _guard1122 & _guard1123;
wire _guard1125 = ev00__0state >= 7'd63;
wire _guard1126 = ev00__0state <= 7'd63;
wire _guard1127 = _guard1125 & _guard1126;
wire _guard1128 = ev00__0state >= 7'd31;
wire _guard1129 = ev00__0state <= 7'd31;
wire _guard1130 = _guard1128 & _guard1129;
wire _guard1131 = ev00__0state >= 7'd95;
wire _guard1132 = ev00__0state <= 7'd95;
wire _guard1133 = _guard1131 & _guard1132;
wire _guard1134 = ev00__0state >= 7'd127;
wire _guard1135 = ev00__0state <= 7'd127;
wire _guard1136 = _guard1134 & _guard1135;
wire _guard1137 = ev00__0state >= 7'd63;
wire _guard1138 = ev00__0state <= 7'd63;
wire _guard1139 = _guard1137 & _guard1138;
wire _guard1140 = ev00__0state >= 7'd31;
wire _guard1141 = ev00__0state <= 7'd31;
wire _guard1142 = _guard1140 & _guard1141;
wire _guard1143 = ev00__0state >= 7'd95;
wire _guard1144 = ev00__0state <= 7'd95;
wire _guard1145 = _guard1143 & _guard1144;
wire _guard1146 = ev00__0state >= 7'd127;
wire _guard1147 = ev00__0state <= 7'd127;
wire _guard1148 = _guard1146 & _guard1147;
wire _guard1149 = ev00__0state >= 7'd63;
wire _guard1150 = ev00__0state <= 7'd63;
wire _guard1151 = _guard1149 & _guard1150;
wire _guard1152 = ev00__0state >= 7'd31;
wire _guard1153 = ev00__0state <= 7'd31;
wire _guard1154 = _guard1152 & _guard1153;
wire _guard1155 = ev00__0state >= 7'd95;
wire _guard1156 = ev00__0state <= 7'd95;
wire _guard1157 = _guard1155 & _guard1156;
wire _guard1158 = ev00__0state >= 7'd127;
wire _guard1159 = ev00__0state <= 7'd127;
wire _guard1160 = _guard1158 & _guard1159;
wire _guard1161 = ev00__0state >= 7'd63;
wire _guard1162 = ev00__0state <= 7'd63;
wire _guard1163 = _guard1161 & _guard1162;
wire _guard1164 = ev00__0state >= 7'd31;
wire _guard1165 = ev00__0state <= 7'd31;
wire _guard1166 = _guard1164 & _guard1165;
wire _guard1167 = ev00__0state >= 7'd95;
wire _guard1168 = ev00__0state <= 7'd95;
wire _guard1169 = _guard1167 & _guard1168;
wire _guard1170 = ev00__0state >= 7'd127;
wire _guard1171 = ev00__0state <= 7'd127;
wire _guard1172 = _guard1170 & _guard1171;
wire _guard1173 = ev00__0state >= 7'd63;
wire _guard1174 = ev00__0state <= 7'd63;
wire _guard1175 = _guard1173 & _guard1174;
wire _guard1176 = ev00__0state >= 7'd31;
wire _guard1177 = ev00__0state <= 7'd31;
wire _guard1178 = _guard1176 & _guard1177;
wire _guard1179 = ev00__0state >= 7'd95;
wire _guard1180 = ev00__0state <= 7'd95;
wire _guard1181 = _guard1179 & _guard1180;
wire _guard1182 = ev00__0state >= 7'd127;
wire _guard1183 = ev00__0state <= 7'd127;
wire _guard1184 = _guard1182 & _guard1183;
wire _guard1185 = ev00__0state >= 7'd63;
wire _guard1186 = ev00__0state <= 7'd63;
wire _guard1187 = _guard1185 & _guard1186;
wire _guard1188 = ev00__0state >= 7'd31;
wire _guard1189 = ev00__0state <= 7'd31;
wire _guard1190 = _guard1188 & _guard1189;
wire _guard1191 = ev00__0state >= 7'd95;
wire _guard1192 = ev00__0state <= 7'd95;
wire _guard1193 = _guard1191 & _guard1192;
wire _guard1194 = ev00__0state >= 7'd127;
wire _guard1195 = ev00__0state <= 7'd127;
wire _guard1196 = _guard1194 & _guard1195;
wire _guard1197 = ev00__0state >= 7'd63;
wire _guard1198 = ev00__0state <= 7'd63;
wire _guard1199 = _guard1197 & _guard1198;
wire _guard1200 = ev00__0state >= 7'd31;
wire _guard1201 = ev00__0state <= 7'd31;
wire _guard1202 = _guard1200 & _guard1201;
wire _guard1203 = ev00__0state >= 7'd95;
wire _guard1204 = ev00__0state <= 7'd95;
wire _guard1205 = _guard1203 & _guard1204;
wire _guard1206 = ev00__0state >= 7'd127;
wire _guard1207 = ev00__0state <= 7'd127;
wire _guard1208 = _guard1206 & _guard1207;
wire _guard1209 = ev00__0state >= 7'd63;
wire _guard1210 = ev00__0state <= 7'd63;
wire _guard1211 = _guard1209 & _guard1210;
wire _guard1212 = ev00__0state >= 7'd31;
wire _guard1213 = ev00__0state <= 7'd31;
wire _guard1214 = _guard1212 & _guard1213;
wire _guard1215 = ev00__0state >= 7'd95;
wire _guard1216 = ev00__0state <= 7'd95;
wire _guard1217 = _guard1215 & _guard1216;
wire _guard1218 = ev00__0state >= 7'd127;
wire _guard1219 = ev00__0state <= 7'd127;
wire _guard1220 = _guard1218 & _guard1219;
wire _guard1221 = ev00__0state >= 7'd63;
wire _guard1222 = ev00__0state <= 7'd63;
wire _guard1223 = _guard1221 & _guard1222;
wire _guard1224 = ev00__0state >= 7'd31;
wire _guard1225 = ev00__0state <= 7'd31;
wire _guard1226 = _guard1224 & _guard1225;
wire _guard1227 = ev00__0state >= 7'd95;
wire _guard1228 = ev00__0state <= 7'd95;
wire _guard1229 = _guard1227 & _guard1228;
wire _guard1230 = ev00__0state >= 7'd127;
wire _guard1231 = ev00__0state <= 7'd127;
wire _guard1232 = _guard1230 & _guard1231;
wire _guard1233 = ev00__0state >= 7'd63;
wire _guard1234 = ev00__0state <= 7'd63;
wire _guard1235 = _guard1233 & _guard1234;
wire _guard1236 = ev00__0state >= 7'd31;
wire _guard1237 = ev00__0state <= 7'd31;
wire _guard1238 = _guard1236 & _guard1237;
wire _guard1239 = ev00__0state >= 7'd95;
wire _guard1240 = ev00__0state <= 7'd95;
wire _guard1241 = _guard1239 & _guard1240;
wire _guard1242 = ev00__0state >= 7'd127;
wire _guard1243 = ev00__0state <= 7'd127;
wire _guard1244 = _guard1242 & _guard1243;
wire _guard1245 = ev00__0state >= 7'd63;
wire _guard1246 = ev00__0state <= 7'd63;
wire _guard1247 = _guard1245 & _guard1246;
wire _guard1248 = ev00__0state >= 7'd31;
wire _guard1249 = ev00__0state <= 7'd31;
wire _guard1250 = _guard1248 & _guard1249;
wire _guard1251 = ev00__0state >= 7'd95;
wire _guard1252 = ev00__0state <= 7'd95;
wire _guard1253 = _guard1251 & _guard1252;
wire _guard1254 = ev00__0state >= 7'd127;
wire _guard1255 = ev00__0state <= 7'd127;
wire _guard1256 = _guard1254 & _guard1255;
wire _guard1257 = ev00__0state >= 7'd63;
wire _guard1258 = ev00__0state <= 7'd63;
wire _guard1259 = _guard1257 & _guard1258;
wire _guard1260 = ev00__0state >= 7'd31;
wire _guard1261 = ev00__0state <= 7'd31;
wire _guard1262 = _guard1260 & _guard1261;
wire _guard1263 = ev00__0state >= 7'd95;
wire _guard1264 = ev00__0state <= 7'd95;
wire _guard1265 = _guard1263 & _guard1264;
wire _guard1266 = ev00__0state >= 7'd127;
wire _guard1267 = ev00__0state <= 7'd127;
wire _guard1268 = _guard1266 & _guard1267;
wire _guard1269 = ev00__0state >= 7'd63;
wire _guard1270 = ev00__0state <= 7'd63;
wire _guard1271 = _guard1269 & _guard1270;
wire _guard1272 = ev00__0state >= 7'd31;
wire _guard1273 = ev00__0state <= 7'd31;
wire _guard1274 = _guard1272 & _guard1273;
wire _guard1275 = ev00__0state >= 7'd95;
wire _guard1276 = ev00__0state <= 7'd95;
wire _guard1277 = _guard1275 & _guard1276;
wire _guard1278 = ev00__0state >= 7'd127;
wire _guard1279 = ev00__0state <= 7'd127;
wire _guard1280 = _guard1278 & _guard1279;
wire _guard1281 = ev00__0state >= 7'd63;
wire _guard1282 = ev00__0state <= 7'd63;
wire _guard1283 = _guard1281 & _guard1282;
wire _guard1284 = ev00__0state >= 7'd31;
wire _guard1285 = ev00__0state <= 7'd31;
wire _guard1286 = _guard1284 & _guard1285;
wire _guard1287 = ev00__0state >= 7'd95;
wire _guard1288 = ev00__0state <= 7'd95;
wire _guard1289 = _guard1287 & _guard1288;
wire _guard1290 = ev00__0state >= 7'd127;
wire _guard1291 = ev00__0state <= 7'd127;
wire _guard1292 = _guard1290 & _guard1291;
wire _guard1293 = ev00__0state >= 7'd63;
wire _guard1294 = ev00__0state <= 7'd63;
wire _guard1295 = _guard1293 & _guard1294;
wire _guard1296 = ev00__0state >= 7'd31;
wire _guard1297 = ev00__0state <= 7'd31;
wire _guard1298 = _guard1296 & _guard1297;
wire _guard1299 = ev00__0state >= 7'd95;
wire _guard1300 = ev00__0state <= 7'd95;
wire _guard1301 = _guard1299 & _guard1300;
wire _guard1302 = ev00__0state >= 7'd127;
wire _guard1303 = ev00__0state <= 7'd127;
wire _guard1304 = _guard1302 & _guard1303;
wire _guard1305 = ev00__0state >= 7'd63;
wire _guard1306 = ev00__0state <= 7'd63;
wire _guard1307 = _guard1305 & _guard1306;
wire _guard1308 = ev00__0state >= 7'd31;
wire _guard1309 = ev00__0state <= 7'd31;
wire _guard1310 = _guard1308 & _guard1309;
wire _guard1311 = ev00__0state >= 7'd95;
wire _guard1312 = ev00__0state <= 7'd95;
wire _guard1313 = _guard1311 & _guard1312;
wire _guard1314 = ev00__0state >= 7'd127;
wire _guard1315 = ev00__0state <= 7'd127;
wire _guard1316 = _guard1314 & _guard1315;
wire _guard1317 = ev00__0state >= 7'd63;
wire _guard1318 = ev00__0state <= 7'd63;
wire _guard1319 = _guard1317 & _guard1318;
wire _guard1320 = ev00__0state >= 7'd31;
wire _guard1321 = ev00__0state <= 7'd31;
wire _guard1322 = _guard1320 & _guard1321;
wire _guard1323 = ev00__0state >= 7'd95;
wire _guard1324 = ev00__0state <= 7'd95;
wire _guard1325 = _guard1323 & _guard1324;
wire _guard1326 = ev00__0state >= 7'd127;
wire _guard1327 = ev00__0state <= 7'd127;
wire _guard1328 = _guard1326 & _guard1327;
wire _guard1329 = ev00__0state >= 7'd63;
wire _guard1330 = ev00__0state <= 7'd63;
wire _guard1331 = _guard1329 & _guard1330;
wire _guard1332 = ev00__0state >= 7'd31;
wire _guard1333 = ev00__0state <= 7'd31;
wire _guard1334 = _guard1332 & _guard1333;
wire _guard1335 = ev00__0state >= 7'd95;
wire _guard1336 = ev00__0state <= 7'd95;
wire _guard1337 = _guard1335 & _guard1336;
wire _guard1338 = ev00__0state >= 7'd127;
wire _guard1339 = ev00__0state <= 7'd127;
wire _guard1340 = _guard1338 & _guard1339;
wire _guard1341 = ev00__0state >= 7'd63;
wire _guard1342 = ev00__0state <= 7'd63;
wire _guard1343 = _guard1341 & _guard1342;
wire _guard1344 = ev00__0state >= 7'd31;
wire _guard1345 = ev00__0state <= 7'd31;
wire _guard1346 = _guard1344 & _guard1345;
wire _guard1347 = ev00__0state >= 7'd95;
wire _guard1348 = ev00__0state <= 7'd95;
wire _guard1349 = _guard1347 & _guard1348;
wire _guard1350 = ev00__0state >= 7'd127;
wire _guard1351 = ev00__0state <= 7'd127;
wire _guard1352 = _guard1350 & _guard1351;
wire _guard1353 = ev00__0state >= 7'd63;
wire _guard1354 = ev00__0state <= 7'd63;
wire _guard1355 = _guard1353 & _guard1354;
wire _guard1356 = ev00__0state >= 7'd31;
wire _guard1357 = ev00__0state <= 7'd31;
wire _guard1358 = _guard1356 & _guard1357;
wire _guard1359 = ev00__0state >= 7'd95;
wire _guard1360 = ev00__0state <= 7'd95;
wire _guard1361 = _guard1359 & _guard1360;
wire _guard1362 = ev00__0state >= 7'd127;
wire _guard1363 = ev00__0state <= 7'd127;
wire _guard1364 = _guard1362 & _guard1363;
wire _guard1365 = ev00__0state >= 7'd63;
wire _guard1366 = ev00__0state <= 7'd63;
wire _guard1367 = _guard1365 & _guard1366;
wire _guard1368 = ev00__0state >= 7'd31;
wire _guard1369 = ev00__0state <= 7'd31;
wire _guard1370 = _guard1368 & _guard1369;
wire _guard1371 = ev00__0state >= 7'd95;
wire _guard1372 = ev00__0state <= 7'd95;
wire _guard1373 = _guard1371 & _guard1372;
wire _guard1374 = ev00__0state >= 7'd127;
wire _guard1375 = ev00__0state <= 7'd127;
wire _guard1376 = _guard1374 & _guard1375;
wire _guard1377 = ev00__0state >= 7'd63;
wire _guard1378 = ev00__0state <= 7'd63;
wire _guard1379 = _guard1377 & _guard1378;
wire _guard1380 = ev00__0state >= 7'd31;
wire _guard1381 = ev00__0state <= 7'd31;
wire _guard1382 = _guard1380 & _guard1381;
wire _guard1383 = ev00__0state >= 7'd95;
wire _guard1384 = ev00__0state <= 7'd95;
wire _guard1385 = _guard1383 & _guard1384;
wire _guard1386 = ev00__0state >= 7'd127;
wire _guard1387 = ev00__0state <= 7'd127;
wire _guard1388 = _guard1386 & _guard1387;
wire _guard1389 = ev00__0state >= 7'd63;
wire _guard1390 = ev00__0state <= 7'd63;
wire _guard1391 = _guard1389 & _guard1390;
wire _guard1392 = ev00__0state >= 7'd31;
wire _guard1393 = ev00__0state <= 7'd31;
wire _guard1394 = _guard1392 & _guard1393;
wire _guard1395 = ev00__0state >= 7'd95;
wire _guard1396 = ev00__0state <= 7'd95;
wire _guard1397 = _guard1395 & _guard1396;
wire _guard1398 = ev00__0state >= 7'd127;
wire _guard1399 = ev00__0state <= 7'd127;
wire _guard1400 = _guard1398 & _guard1399;
wire _guard1401 = ev00__0state >= 7'd63;
wire _guard1402 = ev00__0state <= 7'd63;
wire _guard1403 = _guard1401 & _guard1402;
wire _guard1404 = ev00__0state >= 7'd31;
wire _guard1405 = ev00__0state <= 7'd31;
wire _guard1406 = _guard1404 & _guard1405;
wire _guard1407 = ev00__0state >= 7'd95;
wire _guard1408 = ev00__0state <= 7'd95;
wire _guard1409 = _guard1407 & _guard1408;
wire _guard1410 = ev00__0state >= 7'd127;
wire _guard1411 = ev00__0state <= 7'd127;
wire _guard1412 = _guard1410 & _guard1411;
wire _guard1413 = ev00__0state >= 7'd63;
wire _guard1414 = ev00__0state <= 7'd63;
wire _guard1415 = _guard1413 & _guard1414;
wire _guard1416 = ev00__0state >= 7'd31;
wire _guard1417 = ev00__0state <= 7'd31;
wire _guard1418 = _guard1416 & _guard1417;
wire _guard1419 = ev00__0state >= 7'd126;
wire _guard1420 = ev00__0state <= 7'd126;
wire _guard1421 = _guard1419 & _guard1420;
wire _guard1422 = ev00__0state >= 7'd126;
wire _guard1423 = ev00__0state <= 7'd126;
wire _guard1424 = _guard1422 & _guard1423;
wire _guard1425 = ev00__0state >= 7'd126;
wire _guard1426 = ev00__0state <= 7'd126;
wire _guard1427 = _guard1425 & _guard1426;
wire _guard1428 = ev00__0state >= 7'd126;
wire _guard1429 = ev00__0state <= 7'd126;
wire _guard1430 = _guard1428 & _guard1429;
wire _guard1431 = ev00__0state >= 7'd126;
wire _guard1432 = ev00__0state <= 7'd126;
wire _guard1433 = _guard1431 & _guard1432;
wire _guard1434 = ev00__0state >= 7'd126;
wire _guard1435 = ev00__0state <= 7'd126;
wire _guard1436 = _guard1434 & _guard1435;
wire _guard1437 = ev00__0state >= 7'd126;
wire _guard1438 = ev00__0state <= 7'd126;
wire _guard1439 = _guard1437 & _guard1438;
wire _guard1440 = ev00__0state >= 7'd126;
wire _guard1441 = ev00__0state <= 7'd126;
wire _guard1442 = _guard1440 & _guard1441;
wire _guard1443 = ev00__0state >= 7'd126;
wire _guard1444 = ev00__0state <= 7'd126;
wire _guard1445 = _guard1443 & _guard1444;
wire _guard1446 = ev00__0state >= 7'd126;
wire _guard1447 = ev00__0state <= 7'd126;
wire _guard1448 = _guard1446 & _guard1447;
wire _guard1449 = ev00__0state >= 7'd126;
wire _guard1450 = ev00__0state <= 7'd126;
wire _guard1451 = _guard1449 & _guard1450;
wire _guard1452 = ev00__0state >= 7'd126;
wire _guard1453 = ev00__0state <= 7'd126;
wire _guard1454 = _guard1452 & _guard1453;
wire _guard1455 = ev00__0state >= 7'd126;
wire _guard1456 = ev00__0state <= 7'd126;
wire _guard1457 = _guard1455 & _guard1456;
wire _guard1458 = ev00__0state >= 7'd126;
wire _guard1459 = ev00__0state <= 7'd126;
wire _guard1460 = _guard1458 & _guard1459;
wire _guard1461 = ev00__0state >= 7'd126;
wire _guard1462 = ev00__0state <= 7'd126;
wire _guard1463 = _guard1461 & _guard1462;
wire _guard1464 = ev00__0state >= 7'd126;
wire _guard1465 = ev00__0state <= 7'd126;
wire _guard1466 = _guard1464 & _guard1465;
wire _guard1467 = ev00__0state >= 7'd126;
wire _guard1468 = ev00__0state <= 7'd126;
wire _guard1469 = _guard1467 & _guard1468;
wire _guard1470 = ev00__0state >= 7'd126;
wire _guard1471 = ev00__0state <= 7'd126;
wire _guard1472 = _guard1470 & _guard1471;
wire _guard1473 = ev00__0state >= 7'd126;
wire _guard1474 = ev00__0state <= 7'd126;
wire _guard1475 = _guard1473 & _guard1474;
wire _guard1476 = ev00__0state >= 7'd126;
wire _guard1477 = ev00__0state <= 7'd126;
wire _guard1478 = _guard1476 & _guard1477;
wire _guard1479 = ev00__0state >= 7'd126;
wire _guard1480 = ev00__0state <= 7'd126;
wire _guard1481 = _guard1479 & _guard1480;
wire _guard1482 = ev00__0state >= 7'd126;
wire _guard1483 = ev00__0state <= 7'd126;
wire _guard1484 = _guard1482 & _guard1483;
wire _guard1485 = ev00__0state >= 7'd126;
wire _guard1486 = ev00__0state <= 7'd126;
wire _guard1487 = _guard1485 & _guard1486;
wire _guard1488 = ev00__0state >= 7'd126;
wire _guard1489 = ev00__0state <= 7'd126;
wire _guard1490 = _guard1488 & _guard1489;
wire _guard1491 = ev00__0state >= 7'd126;
wire _guard1492 = ev00__0state <= 7'd126;
wire _guard1493 = _guard1491 & _guard1492;
wire _guard1494 = ev00__0state >= 7'd126;
wire _guard1495 = ev00__0state <= 7'd126;
wire _guard1496 = _guard1494 & _guard1495;
wire _guard1497 = ev00__0state >= 7'd126;
wire _guard1498 = ev00__0state <= 7'd126;
wire _guard1499 = _guard1497 & _guard1498;
wire _guard1500 = ev00__0state >= 7'd126;
wire _guard1501 = ev00__0state <= 7'd126;
wire _guard1502 = _guard1500 & _guard1501;
wire _guard1503 = ev00__0state >= 7'd126;
wire _guard1504 = ev00__0state <= 7'd126;
wire _guard1505 = _guard1503 & _guard1504;
wire _guard1506 = ev00__0state >= 7'd126;
wire _guard1507 = ev00__0state <= 7'd126;
wire _guard1508 = _guard1506 & _guard1507;
wire _guard1509 = ev00__0state >= 7'd126;
wire _guard1510 = ev00__0state <= 7'd126;
wire _guard1511 = _guard1509 & _guard1510;
wire _guard1512 = ev00__0state >= 7'd126;
wire _guard1513 = ev00__0state <= 7'd126;
wire _guard1514 = _guard1512 & _guard1513;
wire _guard1515 = ev00__0state >= 7'd32;
wire _guard1516 = ev00__0state <= 7'd32;
wire _guard1517 = _guard1515 & _guard1516;
wire _guard1518 = ev00__0state >= 7'd64;
wire _guard1519 = ev00__0state <= 7'd64;
wire _guard1520 = _guard1518 & _guard1519;
wire _guard1521 = ev00__0state >= 7'd96;
wire _guard1522 = ev00__0state <= 7'd96;
wire _guard1523 = _guard1521 & _guard1522;
wire _guard1524 = ev00__0_0;
wire _guard1525 = ev00__0state >= 7'd1;
wire _guard1526 = ev00__0state <= 7'd0;
wire _guard1527 = _guard1525 & _guard1526;
wire _guard1528 = _guard1524 | _guard1527;
wire _guard1529 = ev00__0state >= 7'd32;
wire _guard1530 = ev00__0state <= 7'd32;
wire _guard1531 = _guard1529 & _guard1530;
wire _guard1532 = ev00__0state >= 7'd64;
wire _guard1533 = ev00__0state <= 7'd64;
wire _guard1534 = _guard1532 & _guard1533;
wire _guard1535 = ev00__0state >= 7'd96;
wire _guard1536 = ev00__0state <= 7'd96;
wire _guard1537 = _guard1535 & _guard1536;
wire _guard1538 = ev00__0_0;
wire _guard1539 = ev00__0state >= 7'd1;
wire _guard1540 = ev00__0state <= 7'd0;
wire _guard1541 = _guard1539 & _guard1540;
wire _guard1542 = _guard1538 | _guard1541;
wire _guard1543 = ev00__0_0;
wire _guard1544 = ev00__0state >= 7'd1;
wire _guard1545 = ev00__0state <= 7'd0;
wire _guard1546 = _guard1544 & _guard1545;
wire _guard1547 = _guard1543 | _guard1546;
wire _guard1548 = ev00__0state >= 7'd96;
wire _guard1549 = ev00__0state <= 7'd96;
wire _guard1550 = _guard1548 & _guard1549;
wire _guard1551 = ev00__0state >= 7'd64;
wire _guard1552 = ev00__0state <= 7'd64;
wire _guard1553 = _guard1551 & _guard1552;
wire _guard1554 = ev00__0state >= 7'd32;
wire _guard1555 = ev00__0state <= 7'd32;
wire _guard1556 = _guard1554 & _guard1555;
wire _guard1557 = ev00__0state >= 7'd32;
wire _guard1558 = ev00__0state <= 7'd32;
wire _guard1559 = _guard1557 & _guard1558;
wire _guard1560 = ev00__0state >= 7'd64;
wire _guard1561 = ev00__0state <= 7'd64;
wire _guard1562 = _guard1560 & _guard1561;
wire _guard1563 = ev00__0state >= 7'd96;
wire _guard1564 = ev00__0state <= 7'd96;
wire _guard1565 = _guard1563 & _guard1564;
wire _guard1566 = ev00__0_0;
wire _guard1567 = ev00__0state >= 7'd1;
wire _guard1568 = ev00__0state <= 7'd0;
wire _guard1569 = _guard1567 & _guard1568;
wire _guard1570 = _guard1566 | _guard1569;
wire _guard1571 = ev00__0state >= 7'd32;
wire _guard1572 = ev00__0state <= 7'd32;
wire _guard1573 = _guard1571 & _guard1572;
wire _guard1574 = ev00__0state >= 7'd64;
wire _guard1575 = ev00__0state <= 7'd64;
wire _guard1576 = _guard1574 & _guard1575;
wire _guard1577 = ev00__0state >= 7'd96;
wire _guard1578 = ev00__0state <= 7'd96;
wire _guard1579 = _guard1577 & _guard1578;
wire _guard1580 = ev00__0_0;
wire _guard1581 = ev00__0state >= 7'd1;
wire _guard1582 = ev00__0state <= 7'd0;
wire _guard1583 = _guard1581 & _guard1582;
wire _guard1584 = _guard1580 | _guard1583;
wire _guard1585 = ev00__0_0;
wire _guard1586 = ev00__0state >= 7'd1;
wire _guard1587 = ev00__0state <= 7'd0;
wire _guard1588 = _guard1586 & _guard1587;
wire _guard1589 = _guard1585 | _guard1588;
wire _guard1590 = ev00__0state >= 7'd32;
wire _guard1591 = ev00__0state <= 7'd32;
wire _guard1592 = _guard1590 & _guard1591;
wire _guard1593 = _guard1589 | _guard1592;
wire _guard1594 = ev00__0state >= 7'd64;
wire _guard1595 = ev00__0state <= 7'd64;
wire _guard1596 = _guard1594 & _guard1595;
wire _guard1597 = _guard1593 | _guard1596;
wire _guard1598 = ev00__0state >= 7'd96;
wire _guard1599 = ev00__0state <= 7'd96;
wire _guard1600 = _guard1598 & _guard1599;
wire _guard1601 = _guard1597 | _guard1600;
wire _guard1602 = ev00__0state >= 7'd32;
wire _guard1603 = ev00__0state <= 7'd32;
wire _guard1604 = _guard1602 & _guard1603;
wire _guard1605 = ev00__0state >= 7'd64;
wire _guard1606 = ev00__0state <= 7'd64;
wire _guard1607 = _guard1605 & _guard1606;
wire _guard1608 = ev00__0state >= 7'd96;
wire _guard1609 = ev00__0state <= 7'd96;
wire _guard1610 = _guard1608 & _guard1609;
wire _guard1611 = ev00__0_0;
wire _guard1612 = ev00__0state >= 7'd1;
wire _guard1613 = ev00__0state <= 7'd0;
wire _guard1614 = _guard1612 & _guard1613;
wire _guard1615 = _guard1611 | _guard1614;
wire _guard1616 = ev00__0state >= 7'd32;
wire _guard1617 = ev00__0state <= 7'd32;
wire _guard1618 = _guard1616 & _guard1617;
wire _guard1619 = ev00__0state >= 7'd64;
wire _guard1620 = ev00__0state <= 7'd64;
wire _guard1621 = _guard1619 & _guard1620;
wire _guard1622 = ev00__0state >= 7'd96;
wire _guard1623 = ev00__0state <= 7'd96;
wire _guard1624 = _guard1622 & _guard1623;
wire _guard1625 = ev00__0_0;
wire _guard1626 = ev00__0state >= 7'd1;
wire _guard1627 = ev00__0state <= 7'd0;
wire _guard1628 = _guard1626 & _guard1627;
wire _guard1629 = _guard1625 | _guard1628;
wire _guard1630 = ev00__0state >= 7'd32;
wire _guard1631 = ev00__0state <= 7'd32;
wire _guard1632 = _guard1630 & _guard1631;
wire _guard1633 = ev00__0state >= 7'd64;
wire _guard1634 = ev00__0state <= 7'd64;
wire _guard1635 = _guard1633 & _guard1634;
wire _guard1636 = ev00__0state >= 7'd96;
wire _guard1637 = ev00__0state <= 7'd96;
wire _guard1638 = _guard1636 & _guard1637;
wire _guard1639 = ev00__0_0;
wire _guard1640 = ev00__0state >= 7'd1;
wire _guard1641 = ev00__0state <= 7'd0;
wire _guard1642 = _guard1640 & _guard1641;
wire _guard1643 = _guard1639 | _guard1642;
wire _guard1644 = ev00__0state >= 7'd32;
wire _guard1645 = ev00__0state <= 7'd32;
wire _guard1646 = _guard1644 & _guard1645;
wire _guard1647 = ev00__0state >= 7'd64;
wire _guard1648 = ev00__0state <= 7'd64;
wire _guard1649 = _guard1647 & _guard1648;
wire _guard1650 = ev00__0state >= 7'd96;
wire _guard1651 = ev00__0state <= 7'd96;
wire _guard1652 = _guard1650 & _guard1651;
wire _guard1653 = ev00__0_0;
wire _guard1654 = ev00__0state >= 7'd1;
wire _guard1655 = ev00__0state <= 7'd0;
wire _guard1656 = _guard1654 & _guard1655;
wire _guard1657 = _guard1653 | _guard1656;
wire _guard1658 = ev00__0_0;
wire _guard1659 = ev00__0state >= 7'd1;
wire _guard1660 = ev00__0state <= 7'd0;
wire _guard1661 = _guard1659 & _guard1660;
wire _guard1662 = _guard1658 | _guard1661;
wire _guard1663 = ev00__0state >= 7'd96;
wire _guard1664 = ev00__0state <= 7'd96;
wire _guard1665 = _guard1663 & _guard1664;
wire _guard1666 = ev00__0state >= 7'd64;
wire _guard1667 = ev00__0state <= 7'd64;
wire _guard1668 = _guard1666 & _guard1667;
wire _guard1669 = ev00__0state >= 7'd32;
wire _guard1670 = ev00__0state <= 7'd32;
wire _guard1671 = _guard1669 & _guard1670;
wire _guard1672 = ev00__0state >= 7'd32;
wire _guard1673 = ev00__0state <= 7'd32;
wire _guard1674 = _guard1672 & _guard1673;
wire _guard1675 = ev00__0state >= 7'd64;
wire _guard1676 = ev00__0state <= 7'd64;
wire _guard1677 = _guard1675 & _guard1676;
wire _guard1678 = ev00__0state >= 7'd96;
wire _guard1679 = ev00__0state <= 7'd96;
wire _guard1680 = _guard1678 & _guard1679;
wire _guard1681 = ev00__0_0;
wire _guard1682 = ev00__0state >= 7'd1;
wire _guard1683 = ev00__0state <= 7'd0;
wire _guard1684 = _guard1682 & _guard1683;
wire _guard1685 = _guard1681 | _guard1684;
wire _guard1686 = ev00__0state >= 7'd32;
wire _guard1687 = ev00__0state <= 7'd32;
wire _guard1688 = _guard1686 & _guard1687;
wire _guard1689 = ev00__0state >= 7'd64;
wire _guard1690 = ev00__0state <= 7'd64;
wire _guard1691 = _guard1689 & _guard1690;
wire _guard1692 = ev00__0state >= 7'd96;
wire _guard1693 = ev00__0state <= 7'd96;
wire _guard1694 = _guard1692 & _guard1693;
wire _guard1695 = ev00__0_0;
wire _guard1696 = ev00__0state >= 7'd1;
wire _guard1697 = ev00__0state <= 7'd0;
wire _guard1698 = _guard1696 & _guard1697;
wire _guard1699 = _guard1695 | _guard1698;
wire _guard1700 = ev00__0state >= 7'd32;
wire _guard1701 = ev00__0state <= 7'd32;
wire _guard1702 = _guard1700 & _guard1701;
wire _guard1703 = ev00__0state >= 7'd64;
wire _guard1704 = ev00__0state <= 7'd64;
wire _guard1705 = _guard1703 & _guard1704;
wire _guard1706 = ev00__0state >= 7'd96;
wire _guard1707 = ev00__0state <= 7'd96;
wire _guard1708 = _guard1706 & _guard1707;
wire _guard1709 = ev00__0_0;
wire _guard1710 = ev00__0state >= 7'd1;
wire _guard1711 = ev00__0state <= 7'd0;
wire _guard1712 = _guard1710 & _guard1711;
wire _guard1713 = _guard1709 | _guard1712;
wire _guard1714 = ev00__0state >= 7'd32;
wire _guard1715 = ev00__0state <= 7'd32;
wire _guard1716 = _guard1714 & _guard1715;
wire _guard1717 = ev00__0state >= 7'd64;
wire _guard1718 = ev00__0state <= 7'd64;
wire _guard1719 = _guard1717 & _guard1718;
wire _guard1720 = ev00__0state >= 7'd96;
wire _guard1721 = ev00__0state <= 7'd96;
wire _guard1722 = _guard1720 & _guard1721;
wire _guard1723 = ev00__0_0;
wire _guard1724 = ev00__0state >= 7'd1;
wire _guard1725 = ev00__0state <= 7'd0;
wire _guard1726 = _guard1724 & _guard1725;
wire _guard1727 = _guard1723 | _guard1726;
wire _guard1728 = ev00__0state >= 7'd32;
wire _guard1729 = ev00__0state <= 7'd32;
wire _guard1730 = _guard1728 & _guard1729;
wire _guard1731 = ev00__0state >= 7'd64;
wire _guard1732 = ev00__0state <= 7'd64;
wire _guard1733 = _guard1731 & _guard1732;
wire _guard1734 = ev00__0state >= 7'd96;
wire _guard1735 = ev00__0state <= 7'd96;
wire _guard1736 = _guard1734 & _guard1735;
wire _guard1737 = ev00__0_0;
wire _guard1738 = ev00__0state >= 7'd1;
wire _guard1739 = ev00__0state <= 7'd0;
wire _guard1740 = _guard1738 & _guard1739;
wire _guard1741 = _guard1737 | _guard1740;
wire _guard1742 = ev00__0state >= 7'd32;
wire _guard1743 = ev00__0state <= 7'd32;
wire _guard1744 = _guard1742 & _guard1743;
wire _guard1745 = ev00__0state >= 7'd64;
wire _guard1746 = ev00__0state <= 7'd64;
wire _guard1747 = _guard1745 & _guard1746;
wire _guard1748 = ev00__0state >= 7'd96;
wire _guard1749 = ev00__0state <= 7'd96;
wire _guard1750 = _guard1748 & _guard1749;
wire _guard1751 = ev00__0_0;
wire _guard1752 = ev00__0state >= 7'd1;
wire _guard1753 = ev00__0state <= 7'd0;
wire _guard1754 = _guard1752 & _guard1753;
wire _guard1755 = _guard1751 | _guard1754;
wire _guard1756 = ev00__0_0;
wire _guard1757 = ev00__0state >= 7'd1;
wire _guard1758 = ev00__0state <= 7'd0;
wire _guard1759 = _guard1757 & _guard1758;
wire _guard1760 = _guard1756 | _guard1759;
wire _guard1761 = ev00__0state >= 7'd96;
wire _guard1762 = ev00__0state <= 7'd96;
wire _guard1763 = _guard1761 & _guard1762;
wire _guard1764 = ev00__0state >= 7'd64;
wire _guard1765 = ev00__0state <= 7'd64;
wire _guard1766 = _guard1764 & _guard1765;
wire _guard1767 = ev00__0state >= 7'd32;
wire _guard1768 = ev00__0state <= 7'd32;
wire _guard1769 = _guard1767 & _guard1768;
wire _guard1770 = ev00__0_0;
wire _guard1771 = ev00__0state >= 7'd1;
wire _guard1772 = ev00__0state <= 7'd0;
wire _guard1773 = _guard1771 & _guard1772;
wire _guard1774 = _guard1770 | _guard1773;
wire _guard1775 = ev00__0state >= 7'd96;
wire _guard1776 = ev00__0state <= 7'd96;
wire _guard1777 = _guard1775 & _guard1776;
wire _guard1778 = ev00__0state >= 7'd64;
wire _guard1779 = ev00__0state <= 7'd64;
wire _guard1780 = _guard1778 & _guard1779;
wire _guard1781 = ev00__0state >= 7'd32;
wire _guard1782 = ev00__0state <= 7'd32;
wire _guard1783 = _guard1781 & _guard1782;
wire _guard1784 = ev00__0state >= 7'd32;
wire _guard1785 = ev00__0state <= 7'd32;
wire _guard1786 = _guard1784 & _guard1785;
wire _guard1787 = ev00__0state >= 7'd64;
wire _guard1788 = ev00__0state <= 7'd64;
wire _guard1789 = _guard1787 & _guard1788;
wire _guard1790 = ev00__0state >= 7'd96;
wire _guard1791 = ev00__0state <= 7'd96;
wire _guard1792 = _guard1790 & _guard1791;
wire _guard1793 = ev00__0_0;
wire _guard1794 = ev00__0state >= 7'd1;
wire _guard1795 = ev00__0state <= 7'd0;
wire _guard1796 = _guard1794 & _guard1795;
wire _guard1797 = _guard1793 | _guard1796;
wire _guard1798 = ev00__0state >= 7'd32;
wire _guard1799 = ev00__0state <= 7'd32;
wire _guard1800 = _guard1798 & _guard1799;
wire _guard1801 = ev00__0state >= 7'd64;
wire _guard1802 = ev00__0state <= 7'd64;
wire _guard1803 = _guard1801 & _guard1802;
wire _guard1804 = ev00__0state >= 7'd96;
wire _guard1805 = ev00__0state <= 7'd96;
wire _guard1806 = _guard1804 & _guard1805;
wire _guard1807 = ev00__0_0;
wire _guard1808 = ev00__0state >= 7'd1;
wire _guard1809 = ev00__0state <= 7'd0;
wire _guard1810 = _guard1808 & _guard1809;
wire _guard1811 = _guard1807 | _guard1810;
wire _guard1812 = ev00__0_0;
wire _guard1813 = ev00__0state >= 7'd1;
wire _guard1814 = ev00__0state <= 7'd0;
wire _guard1815 = _guard1813 & _guard1814;
wire _guard1816 = _guard1812 | _guard1815;
wire _guard1817 = ev00__0state >= 7'd96;
wire _guard1818 = ev00__0state <= 7'd96;
wire _guard1819 = _guard1817 & _guard1818;
wire _guard1820 = ev00__0state >= 7'd64;
wire _guard1821 = ev00__0state <= 7'd64;
wire _guard1822 = _guard1820 & _guard1821;
wire _guard1823 = ev00__0state >= 7'd32;
wire _guard1824 = ev00__0state <= 7'd32;
wire _guard1825 = _guard1823 & _guard1824;
wire _guard1826 = ev00__0state >= 7'd32;
wire _guard1827 = ev00__0state <= 7'd32;
wire _guard1828 = _guard1826 & _guard1827;
wire _guard1829 = ev00__0state >= 7'd64;
wire _guard1830 = ev00__0state <= 7'd64;
wire _guard1831 = _guard1829 & _guard1830;
wire _guard1832 = ev00__0state >= 7'd96;
wire _guard1833 = ev00__0state <= 7'd96;
wire _guard1834 = _guard1832 & _guard1833;
wire _guard1835 = ev00__0_0;
wire _guard1836 = ev00__0state >= 7'd1;
wire _guard1837 = ev00__0state <= 7'd0;
wire _guard1838 = _guard1836 & _guard1837;
wire _guard1839 = _guard1835 | _guard1838;
wire _guard1840 = ev00__0state >= 7'd32;
wire _guard1841 = ev00__0state <= 7'd32;
wire _guard1842 = _guard1840 & _guard1841;
wire _guard1843 = ev00__0state >= 7'd64;
wire _guard1844 = ev00__0state <= 7'd64;
wire _guard1845 = _guard1843 & _guard1844;
wire _guard1846 = ev00__0state >= 7'd96;
wire _guard1847 = ev00__0state <= 7'd96;
wire _guard1848 = _guard1846 & _guard1847;
wire _guard1849 = ev00__0_0;
wire _guard1850 = ev00__0state >= 7'd1;
wire _guard1851 = ev00__0state <= 7'd0;
wire _guard1852 = _guard1850 & _guard1851;
wire _guard1853 = _guard1849 | _guard1852;
wire _guard1854 = ev00__0_0;
wire _guard1855 = ev00__0state >= 7'd1;
wire _guard1856 = ev00__0state <= 7'd0;
wire _guard1857 = _guard1855 & _guard1856;
wire _guard1858 = _guard1854 | _guard1857;
wire _guard1859 = ev00__0state >= 7'd96;
wire _guard1860 = ev00__0state <= 7'd96;
wire _guard1861 = _guard1859 & _guard1860;
wire _guard1862 = ev00__0state >= 7'd64;
wire _guard1863 = ev00__0state <= 7'd64;
wire _guard1864 = _guard1862 & _guard1863;
wire _guard1865 = ev00__0state >= 7'd32;
wire _guard1866 = ev00__0state <= 7'd32;
wire _guard1867 = _guard1865 & _guard1866;
wire _guard1868 = ev00__0_0;
wire _guard1869 = ev00__0state >= 7'd1;
wire _guard1870 = ev00__0state <= 7'd0;
wire _guard1871 = _guard1869 & _guard1870;
wire _guard1872 = _guard1868 | _guard1871;
wire _guard1873 = ev00__0state >= 7'd96;
wire _guard1874 = ev00__0state <= 7'd96;
wire _guard1875 = _guard1873 & _guard1874;
wire _guard1876 = ev00__0state >= 7'd64;
wire _guard1877 = ev00__0state <= 7'd64;
wire _guard1878 = _guard1876 & _guard1877;
wire _guard1879 = ev00__0state >= 7'd32;
wire _guard1880 = ev00__0state <= 7'd32;
wire _guard1881 = _guard1879 & _guard1880;
wire _guard1882 = ev00__0state >= 7'd32;
wire _guard1883 = ev00__0state <= 7'd32;
wire _guard1884 = _guard1882 & _guard1883;
wire _guard1885 = ev00__0state >= 7'd64;
wire _guard1886 = ev00__0state <= 7'd64;
wire _guard1887 = _guard1885 & _guard1886;
wire _guard1888 = ev00__0state >= 7'd96;
wire _guard1889 = ev00__0state <= 7'd96;
wire _guard1890 = _guard1888 & _guard1889;
wire _guard1891 = ev00__0_0;
wire _guard1892 = ev00__0state >= 7'd1;
wire _guard1893 = ev00__0state <= 7'd0;
wire _guard1894 = _guard1892 & _guard1893;
wire _guard1895 = _guard1891 | _guard1894;
wire _guard1896 = ev00__0_0;
wire _guard1897 = ev00__0state >= 7'd1;
wire _guard1898 = ev00__0state <= 7'd0;
wire _guard1899 = _guard1897 & _guard1898;
wire _guard1900 = _guard1896 | _guard1899;
wire _guard1901 = ev00__0state >= 7'd96;
wire _guard1902 = ev00__0state <= 7'd96;
wire _guard1903 = _guard1901 & _guard1902;
wire _guard1904 = ev00__0state >= 7'd64;
wire _guard1905 = ev00__0state <= 7'd64;
wire _guard1906 = _guard1904 & _guard1905;
wire _guard1907 = ev00__0state >= 7'd32;
wire _guard1908 = ev00__0state <= 7'd32;
wire _guard1909 = _guard1907 & _guard1908;
wire _guard1910 = ev00__0state >= 7'd32;
wire _guard1911 = ev00__0state <= 7'd32;
wire _guard1912 = _guard1910 & _guard1911;
wire _guard1913 = ev00__0state >= 7'd64;
wire _guard1914 = ev00__0state <= 7'd64;
wire _guard1915 = _guard1913 & _guard1914;
wire _guard1916 = ev00__0state >= 7'd96;
wire _guard1917 = ev00__0state <= 7'd96;
wire _guard1918 = _guard1916 & _guard1917;
wire _guard1919 = ev00__0_0;
wire _guard1920 = ev00__0state >= 7'd1;
wire _guard1921 = ev00__0state <= 7'd0;
wire _guard1922 = _guard1920 & _guard1921;
wire _guard1923 = _guard1919 | _guard1922;
wire _guard1924 = ev00__0state >= 7'd32;
wire _guard1925 = ev00__0state <= 7'd32;
wire _guard1926 = _guard1924 & _guard1925;
wire _guard1927 = ev00__0state >= 7'd64;
wire _guard1928 = ev00__0state <= 7'd64;
wire _guard1929 = _guard1927 & _guard1928;
wire _guard1930 = ev00__0state >= 7'd96;
wire _guard1931 = ev00__0state <= 7'd96;
wire _guard1932 = _guard1930 & _guard1931;
wire _guard1933 = ev00__0_0;
wire _guard1934 = ev00__0state >= 7'd1;
wire _guard1935 = ev00__0state <= 7'd0;
wire _guard1936 = _guard1934 & _guard1935;
wire _guard1937 = _guard1933 | _guard1936;
wire _guard1938 = ev00__0_0;
wire _guard1939 = ev00__0state >= 7'd1;
wire _guard1940 = ev00__0state <= 7'd0;
wire _guard1941 = _guard1939 & _guard1940;
wire _guard1942 = _guard1938 | _guard1941;
wire _guard1943 = ev00__0state >= 7'd96;
wire _guard1944 = ev00__0state <= 7'd96;
wire _guard1945 = _guard1943 & _guard1944;
wire _guard1946 = ev00__0state >= 7'd64;
wire _guard1947 = ev00__0state <= 7'd64;
wire _guard1948 = _guard1946 & _guard1947;
wire _guard1949 = ev00__0state >= 7'd32;
wire _guard1950 = ev00__0state <= 7'd32;
wire _guard1951 = _guard1949 & _guard1950;
wire _guard1952 = ev00__0state >= 7'd32;
wire _guard1953 = ev00__0state <= 7'd32;
wire _guard1954 = _guard1952 & _guard1953;
wire _guard1955 = ev00__0state >= 7'd64;
wire _guard1956 = ev00__0state <= 7'd64;
wire _guard1957 = _guard1955 & _guard1956;
wire _guard1958 = ev00__0state >= 7'd96;
wire _guard1959 = ev00__0state <= 7'd96;
wire _guard1960 = _guard1958 & _guard1959;
wire _guard1961 = ev00__0_0;
wire _guard1962 = ev00__0state >= 7'd1;
wire _guard1963 = ev00__0state <= 7'd0;
wire _guard1964 = _guard1962 & _guard1963;
wire _guard1965 = _guard1961 | _guard1964;
wire _guard1966 = ev00__0state >= 7'd32;
wire _guard1967 = ev00__0state <= 7'd32;
wire _guard1968 = _guard1966 & _guard1967;
wire _guard1969 = ev00__0state >= 7'd64;
wire _guard1970 = ev00__0state <= 7'd64;
wire _guard1971 = _guard1969 & _guard1970;
wire _guard1972 = ev00__0state >= 7'd96;
wire _guard1973 = ev00__0state <= 7'd96;
wire _guard1974 = _guard1972 & _guard1973;
wire _guard1975 = ev00__0_0;
wire _guard1976 = ev00__0state >= 7'd1;
wire _guard1977 = ev00__0state <= 7'd0;
wire _guard1978 = _guard1976 & _guard1977;
wire _guard1979 = _guard1975 | _guard1978;
wire _guard1980 = ev00__0_0;
wire _guard1981 = ev00__0state >= 7'd1;
wire _guard1982 = ev00__0state <= 7'd0;
wire _guard1983 = _guard1981 & _guard1982;
wire _guard1984 = _guard1980 | _guard1983;
wire _guard1985 = ev00__0state >= 7'd96;
wire _guard1986 = ev00__0state <= 7'd96;
wire _guard1987 = _guard1985 & _guard1986;
wire _guard1988 = ev00__0state >= 7'd64;
wire _guard1989 = ev00__0state <= 7'd64;
wire _guard1990 = _guard1988 & _guard1989;
wire _guard1991 = ev00__0state >= 7'd32;
wire _guard1992 = ev00__0state <= 7'd32;
wire _guard1993 = _guard1991 & _guard1992;
wire _guard1994 = ev00__0_0;
wire _guard1995 = ev00__0state >= 7'd1;
wire _guard1996 = ev00__0state <= 7'd0;
wire _guard1997 = _guard1995 & _guard1996;
wire _guard1998 = _guard1994 | _guard1997;
wire _guard1999 = ev00__0state >= 7'd96;
wire _guard2000 = ev00__0state <= 7'd96;
wire _guard2001 = _guard1999 & _guard2000;
wire _guard2002 = ev00__0state >= 7'd64;
wire _guard2003 = ev00__0state <= 7'd64;
wire _guard2004 = _guard2002 & _guard2003;
wire _guard2005 = ev00__0state >= 7'd32;
wire _guard2006 = ev00__0state <= 7'd32;
wire _guard2007 = _guard2005 & _guard2006;
wire _guard2008 = ev00__0state >= 7'd32;
wire _guard2009 = ev00__0state <= 7'd32;
wire _guard2010 = _guard2008 & _guard2009;
wire _guard2011 = ev00__0state >= 7'd64;
wire _guard2012 = ev00__0state <= 7'd64;
wire _guard2013 = _guard2011 & _guard2012;
wire _guard2014 = ev00__0state >= 7'd96;
wire _guard2015 = ev00__0state <= 7'd96;
wire _guard2016 = _guard2014 & _guard2015;
wire _guard2017 = ev00__0_0;
wire _guard2018 = ev00__0state >= 7'd1;
wire _guard2019 = ev00__0state <= 7'd0;
wire _guard2020 = _guard2018 & _guard2019;
wire _guard2021 = _guard2017 | _guard2020;
wire _guard2022 = ev00__0state >= 7'd32;
wire _guard2023 = ev00__0state <= 7'd32;
wire _guard2024 = _guard2022 & _guard2023;
wire _guard2025 = ev00__0state >= 7'd64;
wire _guard2026 = ev00__0state <= 7'd64;
wire _guard2027 = _guard2025 & _guard2026;
wire _guard2028 = ev00__0state >= 7'd96;
wire _guard2029 = ev00__0state <= 7'd96;
wire _guard2030 = _guard2028 & _guard2029;
wire _guard2031 = ev00__0_0;
wire _guard2032 = ev00__0state >= 7'd1;
wire _guard2033 = ev00__0state <= 7'd0;
wire _guard2034 = _guard2032 & _guard2033;
wire _guard2035 = _guard2031 | _guard2034;
wire _guard2036 = ev00__0state >= 7'd32;
wire _guard2037 = ev00__0state <= 7'd32;
wire _guard2038 = _guard2036 & _guard2037;
wire _guard2039 = ev00__0state >= 7'd64;
wire _guard2040 = ev00__0state <= 7'd64;
wire _guard2041 = _guard2039 & _guard2040;
wire _guard2042 = ev00__0state >= 7'd96;
wire _guard2043 = ev00__0state <= 7'd96;
wire _guard2044 = _guard2042 & _guard2043;
wire _guard2045 = ev00__0_0;
wire _guard2046 = ev00__0state >= 7'd1;
wire _guard2047 = ev00__0state <= 7'd0;
wire _guard2048 = _guard2046 & _guard2047;
wire _guard2049 = _guard2045 | _guard2048;
wire _guard2050 = ev00__0_0;
wire _guard2051 = ev00__0state >= 7'd1;
wire _guard2052 = ev00__0state <= 7'd0;
wire _guard2053 = _guard2051 & _guard2052;
wire _guard2054 = _guard2050 | _guard2053;
wire _guard2055 = ev00__0state >= 7'd96;
wire _guard2056 = ev00__0state <= 7'd96;
wire _guard2057 = _guard2055 & _guard2056;
wire _guard2058 = ev00__0state >= 7'd64;
wire _guard2059 = ev00__0state <= 7'd64;
wire _guard2060 = _guard2058 & _guard2059;
wire _guard2061 = ev00__0state >= 7'd32;
wire _guard2062 = ev00__0state <= 7'd32;
wire _guard2063 = _guard2061 & _guard2062;
wire _guard2064 = ev00__0state >= 7'd32;
wire _guard2065 = ev00__0state <= 7'd32;
wire _guard2066 = _guard2064 & _guard2065;
wire _guard2067 = ev00__0state >= 7'd64;
wire _guard2068 = ev00__0state <= 7'd64;
wire _guard2069 = _guard2067 & _guard2068;
wire _guard2070 = ev00__0state >= 7'd96;
wire _guard2071 = ev00__0state <= 7'd96;
wire _guard2072 = _guard2070 & _guard2071;
wire _guard2073 = ev00__0_0;
wire _guard2074 = ev00__0state >= 7'd1;
wire _guard2075 = ev00__0state <= 7'd0;
wire _guard2076 = _guard2074 & _guard2075;
wire _guard2077 = _guard2073 | _guard2076;
wire _guard2078 = ev00__0state >= 7'd32;
wire _guard2079 = ev00__0state <= 7'd32;
wire _guard2080 = _guard2078 & _guard2079;
wire _guard2081 = ev00__0state >= 7'd64;
wire _guard2082 = ev00__0state <= 7'd64;
wire _guard2083 = _guard2081 & _guard2082;
wire _guard2084 = ev00__0state >= 7'd96;
wire _guard2085 = ev00__0state <= 7'd96;
wire _guard2086 = _guard2084 & _guard2085;
wire _guard2087 = ev00__0_0;
wire _guard2088 = ev00__0state >= 7'd1;
wire _guard2089 = ev00__0state <= 7'd0;
wire _guard2090 = _guard2088 & _guard2089;
wire _guard2091 = _guard2087 | _guard2090;
wire _guard2092 = ev00__0_0;
wire _guard2093 = ev00__0state >= 7'd1;
wire _guard2094 = ev00__0state <= 7'd0;
wire _guard2095 = _guard2093 & _guard2094;
wire _guard2096 = _guard2092 | _guard2095;
wire _guard2097 = ev00__0state >= 7'd96;
wire _guard2098 = ev00__0state <= 7'd96;
wire _guard2099 = _guard2097 & _guard2098;
wire _guard2100 = ev00__0state >= 7'd64;
wire _guard2101 = ev00__0state <= 7'd64;
wire _guard2102 = _guard2100 & _guard2101;
wire _guard2103 = ev00__0state >= 7'd32;
wire _guard2104 = ev00__0state <= 7'd32;
wire _guard2105 = _guard2103 & _guard2104;
wire _guard2106 = ev00__0state >= 7'd32;
wire _guard2107 = ev00__0state <= 7'd32;
wire _guard2108 = _guard2106 & _guard2107;
wire _guard2109 = ev00__0state >= 7'd64;
wire _guard2110 = ev00__0state <= 7'd64;
wire _guard2111 = _guard2109 & _guard2110;
wire _guard2112 = ev00__0state >= 7'd96;
wire _guard2113 = ev00__0state <= 7'd96;
wire _guard2114 = _guard2112 & _guard2113;
wire _guard2115 = ev00__0_0;
wire _guard2116 = ev00__0state >= 7'd1;
wire _guard2117 = ev00__0state <= 7'd0;
wire _guard2118 = _guard2116 & _guard2117;
wire _guard2119 = _guard2115 | _guard2118;
wire _guard2120 = ev00__0_0;
wire _guard2121 = ev00__0state >= 7'd1;
wire _guard2122 = ev00__0state <= 7'd0;
wire _guard2123 = _guard2121 & _guard2122;
wire _guard2124 = _guard2120 | _guard2123;
wire _guard2125 = ev00__0state >= 7'd96;
wire _guard2126 = ev00__0state <= 7'd96;
wire _guard2127 = _guard2125 & _guard2126;
wire _guard2128 = ev00__0state >= 7'd64;
wire _guard2129 = ev00__0state <= 7'd64;
wire _guard2130 = _guard2128 & _guard2129;
wire _guard2131 = ev00__0state >= 7'd32;
wire _guard2132 = ev00__0state <= 7'd32;
wire _guard2133 = _guard2131 & _guard2132;
wire _guard2134 = ev00__0_0;
wire _guard2135 = ev00__0state >= 7'd1;
wire _guard2136 = ev00__0state <= 7'd0;
wire _guard2137 = _guard2135 & _guard2136;
wire _guard2138 = _guard2134 | _guard2137;
wire _guard2139 = ev00__0state >= 7'd96;
wire _guard2140 = ev00__0state <= 7'd96;
wire _guard2141 = _guard2139 & _guard2140;
wire _guard2142 = ev00__0state >= 7'd64;
wire _guard2143 = ev00__0state <= 7'd64;
wire _guard2144 = _guard2142 & _guard2143;
wire _guard2145 = ev00__0state >= 7'd32;
wire _guard2146 = ev00__0state <= 7'd32;
wire _guard2147 = _guard2145 & _guard2146;
wire _guard2148 = ev00__0state >= 7'd32;
wire _guard2149 = ev00__0state <= 7'd32;
wire _guard2150 = _guard2148 & _guard2149;
wire _guard2151 = ev00__0state >= 7'd64;
wire _guard2152 = ev00__0state <= 7'd64;
wire _guard2153 = _guard2151 & _guard2152;
wire _guard2154 = ev00__0state >= 7'd96;
wire _guard2155 = ev00__0state <= 7'd96;
wire _guard2156 = _guard2154 & _guard2155;
wire _guard2157 = ev00__0_0;
wire _guard2158 = ev00__0state >= 7'd1;
wire _guard2159 = ev00__0state <= 7'd0;
wire _guard2160 = _guard2158 & _guard2159;
wire _guard2161 = _guard2157 | _guard2160;
wire _guard2162 = ev00__0state >= 7'd32;
wire _guard2163 = ev00__0state <= 7'd32;
wire _guard2164 = _guard2162 & _guard2163;
wire _guard2165 = ev00__0state >= 7'd64;
wire _guard2166 = ev00__0state <= 7'd64;
wire _guard2167 = _guard2165 & _guard2166;
wire _guard2168 = ev00__0state >= 7'd96;
wire _guard2169 = ev00__0state <= 7'd96;
wire _guard2170 = _guard2168 & _guard2169;
wire _guard2171 = ev00__0_0;
wire _guard2172 = ev00__0state >= 7'd1;
wire _guard2173 = ev00__0state <= 7'd0;
wire _guard2174 = _guard2172 & _guard2173;
wire _guard2175 = _guard2171 | _guard2174;
wire _guard2176 = ev00__0state >= 7'd32;
wire _guard2177 = ev00__0state <= 7'd32;
wire _guard2178 = _guard2176 & _guard2177;
wire _guard2179 = ev00__0state >= 7'd64;
wire _guard2180 = ev00__0state <= 7'd64;
wire _guard2181 = _guard2179 & _guard2180;
wire _guard2182 = ev00__0state >= 7'd96;
wire _guard2183 = ev00__0state <= 7'd96;
wire _guard2184 = _guard2182 & _guard2183;
wire _guard2185 = ev00__0_0;
wire _guard2186 = ev00__0state >= 7'd1;
wire _guard2187 = ev00__0state <= 7'd0;
wire _guard2188 = _guard2186 & _guard2187;
wire _guard2189 = _guard2185 | _guard2188;
wire _guard2190 = ev00__0_0;
wire _guard2191 = ev00__0state >= 7'd1;
wire _guard2192 = ev00__0state <= 7'd0;
wire _guard2193 = _guard2191 & _guard2192;
wire _guard2194 = _guard2190 | _guard2193;
wire _guard2195 = ev00__0state >= 7'd96;
wire _guard2196 = ev00__0state <= 7'd96;
wire _guard2197 = _guard2195 & _guard2196;
wire _guard2198 = ev00__0state >= 7'd64;
wire _guard2199 = ev00__0state <= 7'd64;
wire _guard2200 = _guard2198 & _guard2199;
wire _guard2201 = ev00__0state >= 7'd32;
wire _guard2202 = ev00__0state <= 7'd32;
wire _guard2203 = _guard2201 & _guard2202;
wire _guard2204 = ev00__0_0;
wire _guard2205 = ev00__0state >= 7'd1;
wire _guard2206 = ev00__0state <= 7'd127;
wire _guard2207 = _guard2205 & _guard2206;
wire _guard2208 = _guard2204 | _guard2207;
wire _guard2209 = ev00__0_0;
wire _guard2210 = ev00__0state >= 7'd1;
wire _guard2211 = ev00__0state <= 7'd127;
wire _guard2212 = _guard2210 & _guard2211;
wire _guard2213 = _guard2209 | _guard2212;
wire _guard2214 = ev00__0_0;
wire _guard2215 = ev00__0state >= 7'd1;
wire _guard2216 = ev00__0state <= 7'd127;
wire _guard2217 = _guard2215 & _guard2216;
wire _guard2218 = _guard2214 | _guard2217;
wire _guard2219 = ev00__0_0;
wire _guard2220 = ev00__0state >= 7'd1;
wire _guard2221 = ev00__0state <= 7'd127;
wire _guard2222 = _guard2220 & _guard2221;
wire _guard2223 = _guard2219 | _guard2222;
wire _guard2224 = ev00__0_0;
wire _guard2225 = ev00__0state >= 7'd1;
wire _guard2226 = ev00__0state <= 7'd127;
wire _guard2227 = _guard2225 & _guard2226;
wire _guard2228 = _guard2224 | _guard2227;
wire _guard2229 = ev00__0_0;
wire _guard2230 = ev00__0state >= 7'd1;
wire _guard2231 = ev00__0state <= 7'd127;
wire _guard2232 = _guard2230 & _guard2231;
wire _guard2233 = _guard2229 | _guard2232;
wire _guard2234 = ev00__0_0;
wire _guard2235 = ev00__0state >= 7'd1;
wire _guard2236 = ev00__0state <= 7'd127;
wire _guard2237 = _guard2235 & _guard2236;
wire _guard2238 = _guard2234 | _guard2237;
wire _guard2239 = ev00__0_0;
wire _guard2240 = ev00__0state >= 7'd1;
wire _guard2241 = ev00__0state <= 7'd127;
wire _guard2242 = _guard2240 & _guard2241;
wire _guard2243 = _guard2239 | _guard2242;
wire _guard2244 = ev00__0_0;
wire _guard2245 = ev00__0state >= 7'd1;
wire _guard2246 = ev00__0state <= 7'd127;
wire _guard2247 = _guard2245 & _guard2246;
wire _guard2248 = _guard2244 | _guard2247;
wire _guard2249 = ev00__0_0;
wire _guard2250 = ev00__0state >= 7'd1;
wire _guard2251 = ev00__0state <= 7'd127;
wire _guard2252 = _guard2250 & _guard2251;
wire _guard2253 = _guard2249 | _guard2252;
wire _guard2254 = ev00__0_0;
wire _guard2255 = ev00__0state >= 7'd1;
wire _guard2256 = ev00__0state <= 7'd127;
wire _guard2257 = _guard2255 & _guard2256;
wire _guard2258 = _guard2254 | _guard2257;
wire _guard2259 = ev00__0_0;
wire _guard2260 = ev00__0state >= 7'd1;
wire _guard2261 = ev00__0state <= 7'd127;
wire _guard2262 = _guard2260 & _guard2261;
wire _guard2263 = _guard2259 | _guard2262;
wire _guard2264 = ev00__0_0;
wire _guard2265 = ev00__0state >= 7'd1;
wire _guard2266 = ev00__0state <= 7'd127;
wire _guard2267 = _guard2265 & _guard2266;
wire _guard2268 = _guard2264 | _guard2267;
wire _guard2269 = ev00__0_0;
wire _guard2270 = ev00__0state >= 7'd1;
wire _guard2271 = ev00__0state <= 7'd127;
wire _guard2272 = _guard2270 & _guard2271;
wire _guard2273 = _guard2269 | _guard2272;
wire _guard2274 = ev00__0_0;
wire _guard2275 = ev00__0state >= 7'd1;
wire _guard2276 = ev00__0state <= 7'd127;
wire _guard2277 = _guard2275 & _guard2276;
wire _guard2278 = _guard2274 | _guard2277;
wire _guard2279 = ev00__0_0;
wire _guard2280 = ev00__0state >= 7'd1;
wire _guard2281 = ev00__0state <= 7'd127;
wire _guard2282 = _guard2280 & _guard2281;
wire _guard2283 = _guard2279 | _guard2282;
wire _guard2284 = ev00__0state >= 7'd96;
wire _guard2285 = ev00__0state <= 7'd96;
wire _guard2286 = _guard2284 & _guard2285;
wire _guard2287 = ev00__0state >= 7'd96;
wire _guard2288 = ev00__0state <= 7'd96;
wire _guard2289 = _guard2287 & _guard2288;
wire _guard2290 = ev00__0state >= 7'd96;
wire _guard2291 = ev00__0state <= 7'd96;
wire _guard2292 = _guard2290 & _guard2291;
wire _guard2293 = ev00__0state >= 7'd96;
wire _guard2294 = ev00__0state <= 7'd96;
wire _guard2295 = _guard2293 & _guard2294;
wire _guard2296 = ev00__0state >= 7'd96;
wire _guard2297 = ev00__0state <= 7'd96;
wire _guard2298 = _guard2296 & _guard2297;
wire _guard2299 = ev00__0state >= 7'd96;
wire _guard2300 = ev00__0state <= 7'd96;
wire _guard2301 = _guard2299 & _guard2300;
wire _guard2302 = ev00__0state >= 7'd96;
wire _guard2303 = ev00__0state <= 7'd96;
wire _guard2304 = _guard2302 & _guard2303;
wire _guard2305 = ev00__0state >= 7'd96;
wire _guard2306 = ev00__0state <= 7'd96;
wire _guard2307 = _guard2305 & _guard2306;
wire _guard2308 = ev00__0state >= 7'd96;
wire _guard2309 = ev00__0state <= 7'd96;
wire _guard2310 = _guard2308 & _guard2309;
wire _guard2311 = ev00__0state >= 7'd96;
wire _guard2312 = ev00__0state <= 7'd96;
wire _guard2313 = _guard2311 & _guard2312;
wire _guard2314 = ev00__0state >= 7'd96;
wire _guard2315 = ev00__0state <= 7'd96;
wire _guard2316 = _guard2314 & _guard2315;
wire _guard2317 = ev00__0state >= 7'd96;
wire _guard2318 = ev00__0state <= 7'd96;
wire _guard2319 = _guard2317 & _guard2318;
wire _guard2320 = ev00__0state >= 7'd96;
wire _guard2321 = ev00__0state <= 7'd96;
wire _guard2322 = _guard2320 & _guard2321;
wire _guard2323 = ev00__0state >= 7'd96;
wire _guard2324 = ev00__0state <= 7'd96;
wire _guard2325 = _guard2323 & _guard2324;
wire _guard2326 = ev00__0state >= 7'd96;
wire _guard2327 = ev00__0state <= 7'd96;
wire _guard2328 = _guard2326 & _guard2327;
wire _guard2329 = ev00__0state >= 7'd96;
wire _guard2330 = ev00__0state <= 7'd96;
wire _guard2331 = _guard2329 & _guard2330;
wire _guard2332 = ev00__0state >= 7'd96;
wire _guard2333 = ev00__0state <= 7'd96;
wire _guard2334 = _guard2332 & _guard2333;
wire _guard2335 = ev00__0state >= 7'd96;
wire _guard2336 = ev00__0state <= 7'd96;
wire _guard2337 = _guard2335 & _guard2336;
wire _guard2338 = ev00__0state >= 7'd96;
wire _guard2339 = ev00__0state <= 7'd96;
wire _guard2340 = _guard2338 & _guard2339;
wire _guard2341 = ev00__0state >= 7'd96;
wire _guard2342 = ev00__0state <= 7'd96;
wire _guard2343 = _guard2341 & _guard2342;
wire _guard2344 = ev00__0state >= 7'd96;
wire _guard2345 = ev00__0state <= 7'd96;
wire _guard2346 = _guard2344 & _guard2345;
wire _guard2347 = ev00__0state >= 7'd96;
wire _guard2348 = ev00__0state <= 7'd96;
wire _guard2349 = _guard2347 & _guard2348;
wire _guard2350 = ev00__0state >= 7'd96;
wire _guard2351 = ev00__0state <= 7'd96;
wire _guard2352 = _guard2350 & _guard2351;
wire _guard2353 = ev00__0state >= 7'd96;
wire _guard2354 = ev00__0state <= 7'd96;
wire _guard2355 = _guard2353 & _guard2354;
wire _guard2356 = ev00__0state >= 7'd96;
wire _guard2357 = ev00__0state <= 7'd96;
wire _guard2358 = _guard2356 & _guard2357;
wire _guard2359 = ev00__0state >= 7'd96;
wire _guard2360 = ev00__0state <= 7'd96;
wire _guard2361 = _guard2359 & _guard2360;
wire _guard2362 = ev00__0state >= 7'd96;
wire _guard2363 = ev00__0state <= 7'd96;
wire _guard2364 = _guard2362 & _guard2363;
wire _guard2365 = ev00__0state >= 7'd96;
wire _guard2366 = ev00__0state <= 7'd96;
wire _guard2367 = _guard2365 & _guard2366;
wire _guard2368 = ev00__0state >= 7'd96;
wire _guard2369 = ev00__0state <= 7'd96;
wire _guard2370 = _guard2368 & _guard2369;
wire _guard2371 = ev00__0state >= 7'd96;
wire _guard2372 = ev00__0state <= 7'd96;
wire _guard2373 = _guard2371 & _guard2372;
wire _guard2374 = ev00__0state >= 7'd96;
wire _guard2375 = ev00__0state <= 7'd96;
wire _guard2376 = _guard2374 & _guard2375;
wire _guard2377 = ev00__0state >= 7'd96;
wire _guard2378 = ev00__0state <= 7'd96;
wire _guard2379 = _guard2377 & _guard2378;
wire _guard2380 = ev00__0state >= 7'd32;
wire _guard2381 = ev00__0state <= 7'd32;
wire _guard2382 = _guard2380 & _guard2381;
wire _guard2383 = ev00__0state >= 7'd95;
wire _guard2384 = ev00__0state <= 7'd95;
wire _guard2385 = _guard2383 & _guard2384;
wire _guard2386 = ev00__0state >= 7'd95;
wire _guard2387 = ev00__0state <= 7'd95;
wire _guard2388 = _guard2386 & _guard2387;
wire _guard2389 = ev00__0state >= 7'd95;
wire _guard2390 = ev00__0state <= 7'd95;
wire _guard2391 = _guard2389 & _guard2390;
wire _guard2392 = ev00__0state >= 7'd95;
wire _guard2393 = ev00__0state <= 7'd95;
wire _guard2394 = _guard2392 & _guard2393;
wire _guard2395 = ev00__0state >= 7'd95;
wire _guard2396 = ev00__0state <= 7'd95;
wire _guard2397 = _guard2395 & _guard2396;
wire _guard2398 = ev00__0state >= 7'd95;
wire _guard2399 = ev00__0state <= 7'd95;
wire _guard2400 = _guard2398 & _guard2399;
wire _guard2401 = ev00__0state >= 7'd95;
wire _guard2402 = ev00__0state <= 7'd95;
wire _guard2403 = _guard2401 & _guard2402;
wire _guard2404 = ev00__0state >= 7'd95;
wire _guard2405 = ev00__0state <= 7'd95;
wire _guard2406 = _guard2404 & _guard2405;
wire _guard2407 = ev00__0state >= 7'd95;
wire _guard2408 = ev00__0state <= 7'd95;
wire _guard2409 = _guard2407 & _guard2408;
wire _guard2410 = ev00__0state >= 7'd95;
wire _guard2411 = ev00__0state <= 7'd95;
wire _guard2412 = _guard2410 & _guard2411;
wire _guard2413 = ev00__0state >= 7'd95;
wire _guard2414 = ev00__0state <= 7'd95;
wire _guard2415 = _guard2413 & _guard2414;
wire _guard2416 = ev00__0state >= 7'd95;
wire _guard2417 = ev00__0state <= 7'd95;
wire _guard2418 = _guard2416 & _guard2417;
wire _guard2419 = ev00__0state >= 7'd95;
wire _guard2420 = ev00__0state <= 7'd95;
wire _guard2421 = _guard2419 & _guard2420;
wire _guard2422 = ev00__0state >= 7'd95;
wire _guard2423 = ev00__0state <= 7'd95;
wire _guard2424 = _guard2422 & _guard2423;
wire _guard2425 = ev00__0state >= 7'd95;
wire _guard2426 = ev00__0state <= 7'd95;
wire _guard2427 = _guard2425 & _guard2426;
wire _guard2428 = ev00__0state >= 7'd95;
wire _guard2429 = ev00__0state <= 7'd95;
wire _guard2430 = _guard2428 & _guard2429;
wire _guard2431 = ev00__0state >= 7'd95;
wire _guard2432 = ev00__0state <= 7'd95;
wire _guard2433 = _guard2431 & _guard2432;
wire _guard2434 = ev00__0state >= 7'd95;
wire _guard2435 = ev00__0state <= 7'd95;
wire _guard2436 = _guard2434 & _guard2435;
wire _guard2437 = ev00__0state >= 7'd95;
wire _guard2438 = ev00__0state <= 7'd95;
wire _guard2439 = _guard2437 & _guard2438;
wire _guard2440 = ev00__0state >= 7'd95;
wire _guard2441 = ev00__0state <= 7'd95;
wire _guard2442 = _guard2440 & _guard2441;
wire _guard2443 = ev00__0state >= 7'd95;
wire _guard2444 = ev00__0state <= 7'd95;
wire _guard2445 = _guard2443 & _guard2444;
wire _guard2446 = ev00__0state >= 7'd95;
wire _guard2447 = ev00__0state <= 7'd95;
wire _guard2448 = _guard2446 & _guard2447;
wire _guard2449 = ev00__0state >= 7'd95;
wire _guard2450 = ev00__0state <= 7'd95;
wire _guard2451 = _guard2449 & _guard2450;
wire _guard2452 = ev00__0state >= 7'd95;
wire _guard2453 = ev00__0state <= 7'd95;
wire _guard2454 = _guard2452 & _guard2453;
wire _guard2455 = ev00__0state >= 7'd95;
wire _guard2456 = ev00__0state <= 7'd95;
wire _guard2457 = _guard2455 & _guard2456;
wire _guard2458 = ev00__0state >= 7'd95;
wire _guard2459 = ev00__0state <= 7'd95;
wire _guard2460 = _guard2458 & _guard2459;
wire _guard2461 = ev00__0state >= 7'd95;
wire _guard2462 = ev00__0state <= 7'd95;
wire _guard2463 = _guard2461 & _guard2462;
wire _guard2464 = ev00__0state >= 7'd95;
wire _guard2465 = ev00__0state <= 7'd95;
wire _guard2466 = _guard2464 & _guard2465;
wire _guard2467 = ev00__0state >= 7'd95;
wire _guard2468 = ev00__0state <= 7'd95;
wire _guard2469 = _guard2467 & _guard2468;
wire _guard2470 = ev00__0state >= 7'd95;
wire _guard2471 = ev00__0state <= 7'd95;
wire _guard2472 = _guard2470 & _guard2471;
wire _guard2473 = ev00__0state >= 7'd95;
wire _guard2474 = ev00__0state <= 7'd95;
wire _guard2475 = _guard2473 & _guard2474;
wire _guard2476 = ev00__0state >= 7'd95;
wire _guard2477 = ev00__0state <= 7'd95;
wire _guard2478 = _guard2476 & _guard2477;
wire _guard2479 = ev00__0state >= 7'd64;
wire _guard2480 = ev00__0state <= 7'd64;
wire _guard2481 = _guard2479 & _guard2480;
wire _guard2482 = ev00__0state >= 7'd64;
wire _guard2483 = ev00__0state <= 7'd64;
wire _guard2484 = _guard2482 & _guard2483;
wire _guard2485 = ev00__0state >= 7'd64;
wire _guard2486 = ev00__0state <= 7'd64;
wire _guard2487 = _guard2485 & _guard2486;
wire _guard2488 = ev00__0state >= 7'd64;
wire _guard2489 = ev00__0state <= 7'd64;
wire _guard2490 = _guard2488 & _guard2489;
wire _guard2491 = ev00__0state >= 7'd64;
wire _guard2492 = ev00__0state <= 7'd64;
wire _guard2493 = _guard2491 & _guard2492;
wire _guard2494 = ev00__0state >= 7'd64;
wire _guard2495 = ev00__0state <= 7'd64;
wire _guard2496 = _guard2494 & _guard2495;
wire _guard2497 = ev00__0state >= 7'd64;
wire _guard2498 = ev00__0state <= 7'd64;
wire _guard2499 = _guard2497 & _guard2498;
wire _guard2500 = ev00__0state >= 7'd64;
wire _guard2501 = ev00__0state <= 7'd64;
wire _guard2502 = _guard2500 & _guard2501;
wire _guard2503 = ev00__0state >= 7'd64;
wire _guard2504 = ev00__0state <= 7'd64;
wire _guard2505 = _guard2503 & _guard2504;
wire _guard2506 = ev00__0state >= 7'd64;
wire _guard2507 = ev00__0state <= 7'd64;
wire _guard2508 = _guard2506 & _guard2507;
wire _guard2509 = ev00__0state >= 7'd64;
wire _guard2510 = ev00__0state <= 7'd64;
wire _guard2511 = _guard2509 & _guard2510;
wire _guard2512 = ev00__0state >= 7'd64;
wire _guard2513 = ev00__0state <= 7'd64;
wire _guard2514 = _guard2512 & _guard2513;
wire _guard2515 = ev00__0state >= 7'd64;
wire _guard2516 = ev00__0state <= 7'd64;
wire _guard2517 = _guard2515 & _guard2516;
wire _guard2518 = ev00__0state >= 7'd64;
wire _guard2519 = ev00__0state <= 7'd64;
wire _guard2520 = _guard2518 & _guard2519;
wire _guard2521 = ev00__0state >= 7'd64;
wire _guard2522 = ev00__0state <= 7'd64;
wire _guard2523 = _guard2521 & _guard2522;
wire _guard2524 = ev00__0state >= 7'd64;
wire _guard2525 = ev00__0state <= 7'd64;
wire _guard2526 = _guard2524 & _guard2525;
wire _guard2527 = ev00__0state >= 7'd64;
wire _guard2528 = ev00__0state <= 7'd64;
wire _guard2529 = _guard2527 & _guard2528;
wire _guard2530 = ev00__0state >= 7'd64;
wire _guard2531 = ev00__0state <= 7'd64;
wire _guard2532 = _guard2530 & _guard2531;
wire _guard2533 = ev00__0state >= 7'd64;
wire _guard2534 = ev00__0state <= 7'd64;
wire _guard2535 = _guard2533 & _guard2534;
wire _guard2536 = ev00__0state >= 7'd64;
wire _guard2537 = ev00__0state <= 7'd64;
wire _guard2538 = _guard2536 & _guard2537;
wire _guard2539 = ev00__0state >= 7'd64;
wire _guard2540 = ev00__0state <= 7'd64;
wire _guard2541 = _guard2539 & _guard2540;
wire _guard2542 = ev00__0state >= 7'd64;
wire _guard2543 = ev00__0state <= 7'd64;
wire _guard2544 = _guard2542 & _guard2543;
wire _guard2545 = ev00__0state >= 7'd64;
wire _guard2546 = ev00__0state <= 7'd64;
wire _guard2547 = _guard2545 & _guard2546;
wire _guard2548 = ev00__0state >= 7'd64;
wire _guard2549 = ev00__0state <= 7'd64;
wire _guard2550 = _guard2548 & _guard2549;
wire _guard2551 = ev00__0state >= 7'd64;
wire _guard2552 = ev00__0state <= 7'd64;
wire _guard2553 = _guard2551 & _guard2552;
wire _guard2554 = ev00__0state >= 7'd64;
wire _guard2555 = ev00__0state <= 7'd64;
wire _guard2556 = _guard2554 & _guard2555;
wire _guard2557 = ev00__0state >= 7'd64;
wire _guard2558 = ev00__0state <= 7'd64;
wire _guard2559 = _guard2557 & _guard2558;
wire _guard2560 = ev00__0state >= 7'd64;
wire _guard2561 = ev00__0state <= 7'd64;
wire _guard2562 = _guard2560 & _guard2561;
wire _guard2563 = ev00__0state >= 7'd64;
wire _guard2564 = ev00__0state <= 7'd64;
wire _guard2565 = _guard2563 & _guard2564;
wire _guard2566 = ev00__0state >= 7'd64;
wire _guard2567 = ev00__0state <= 7'd64;
wire _guard2568 = _guard2566 & _guard2567;
wire _guard2569 = ev00__0state >= 7'd64;
wire _guard2570 = ev00__0state <= 7'd64;
wire _guard2571 = _guard2569 & _guard2570;
wire _guard2572 = ev00__0state >= 7'd64;
wire _guard2573 = ev00__0state <= 7'd64;
wire _guard2574 = _guard2572 & _guard2573;
wire _guard2575 = ev00__0_0;
wire _guard2576 = ev00__0state >= 7'd1;
wire _guard2577 = ev00__0state <= 7'd127;
wire _guard2578 = _guard2576 & _guard2577;
wire _guard2579 = _guard2575 | _guard2578;
wire _guard2580 = ev00__0_0;
wire _guard2581 = ev00__0state >= 7'd1;
wire _guard2582 = ev00__0state <= 7'd127;
wire _guard2583 = _guard2581 & _guard2582;
wire _guard2584 = _guard2580 | _guard2583;
wire _guard2585 = ev00__0_0;
wire _guard2586 = ev00__0state >= 7'd1;
wire _guard2587 = ev00__0state <= 7'd127;
wire _guard2588 = _guard2586 & _guard2587;
wire _guard2589 = _guard2585 | _guard2588;
wire _guard2590 = ev00__0_0;
wire _guard2591 = ev00__0state >= 7'd1;
wire _guard2592 = ev00__0state <= 7'd127;
wire _guard2593 = _guard2591 & _guard2592;
wire _guard2594 = _guard2590 | _guard2593;
wire _guard2595 = ev00__0_0;
wire _guard2596 = ev00__0state >= 7'd1;
wire _guard2597 = ev00__0state <= 7'd127;
wire _guard2598 = _guard2596 & _guard2597;
wire _guard2599 = _guard2595 | _guard2598;
wire _guard2600 = ev00__0_0;
wire _guard2601 = ev00__0state >= 7'd1;
wire _guard2602 = ev00__0state <= 7'd127;
wire _guard2603 = _guard2601 & _guard2602;
wire _guard2604 = _guard2600 | _guard2603;
wire _guard2605 = ev00__0_0;
wire _guard2606 = ev00__0state >= 7'd1;
wire _guard2607 = ev00__0state <= 7'd127;
wire _guard2608 = _guard2606 & _guard2607;
wire _guard2609 = _guard2605 | _guard2608;
wire _guard2610 = ev00__0_0;
wire _guard2611 = ev00__0state >= 7'd1;
wire _guard2612 = ev00__0state <= 7'd127;
wire _guard2613 = _guard2611 & _guard2612;
wire _guard2614 = _guard2610 | _guard2613;
wire _guard2615 = ev00__0_0;
wire _guard2616 = ev00__0state >= 7'd1;
wire _guard2617 = ev00__0state <= 7'd127;
wire _guard2618 = _guard2616 & _guard2617;
wire _guard2619 = _guard2615 | _guard2618;
wire _guard2620 = ev00__0_0;
wire _guard2621 = ev00__0state >= 7'd1;
wire _guard2622 = ev00__0state <= 7'd127;
wire _guard2623 = _guard2621 & _guard2622;
wire _guard2624 = _guard2620 | _guard2623;
wire _guard2625 = ev00__0_0;
wire _guard2626 = ev00__0state >= 7'd1;
wire _guard2627 = ev00__0state <= 7'd127;
wire _guard2628 = _guard2626 & _guard2627;
wire _guard2629 = _guard2625 | _guard2628;
wire _guard2630 = ev00__0_0;
wire _guard2631 = ev00__0state >= 7'd1;
wire _guard2632 = ev00__0state <= 7'd127;
wire _guard2633 = _guard2631 & _guard2632;
wire _guard2634 = _guard2630 | _guard2633;
wire _guard2635 = ev00__0_0;
wire _guard2636 = ev00__0state >= 7'd1;
wire _guard2637 = ev00__0state <= 7'd127;
wire _guard2638 = _guard2636 & _guard2637;
wire _guard2639 = _guard2635 | _guard2638;
wire _guard2640 = ev00__0_0;
wire _guard2641 = ev00__0state >= 7'd1;
wire _guard2642 = ev00__0state <= 7'd127;
wire _guard2643 = _guard2641 & _guard2642;
wire _guard2644 = _guard2640 | _guard2643;
wire _guard2645 = ev00__0_0;
wire _guard2646 = ev00__0state >= 7'd1;
wire _guard2647 = ev00__0state <= 7'd127;
wire _guard2648 = _guard2646 & _guard2647;
wire _guard2649 = _guard2645 | _guard2648;
wire _guard2650 = ev00__0_0;
wire _guard2651 = ev00__0state >= 7'd1;
wire _guard2652 = ev00__0state <= 7'd127;
wire _guard2653 = _guard2651 & _guard2652;
wire _guard2654 = _guard2650 | _guard2653;
wire _guard2655 = ev00__0state >= 7'd94;
wire _guard2656 = ev00__0state <= 7'd94;
wire _guard2657 = _guard2655 & _guard2656;
wire _guard2658 = ev00__0state >= 7'd94;
wire _guard2659 = ev00__0state <= 7'd94;
wire _guard2660 = _guard2658 & _guard2659;
wire _guard2661 = ev00__0state >= 7'd94;
wire _guard2662 = ev00__0state <= 7'd94;
wire _guard2663 = _guard2661 & _guard2662;
wire _guard2664 = ev00__0state >= 7'd94;
wire _guard2665 = ev00__0state <= 7'd94;
wire _guard2666 = _guard2664 & _guard2665;
wire _guard2667 = ev00__0state >= 7'd94;
wire _guard2668 = ev00__0state <= 7'd94;
wire _guard2669 = _guard2667 & _guard2668;
wire _guard2670 = ev00__0state >= 7'd94;
wire _guard2671 = ev00__0state <= 7'd94;
wire _guard2672 = _guard2670 & _guard2671;
wire _guard2673 = ev00__0state >= 7'd94;
wire _guard2674 = ev00__0state <= 7'd94;
wire _guard2675 = _guard2673 & _guard2674;
wire _guard2676 = ev00__0state >= 7'd94;
wire _guard2677 = ev00__0state <= 7'd94;
wire _guard2678 = _guard2676 & _guard2677;
wire _guard2679 = ev00__0state >= 7'd94;
wire _guard2680 = ev00__0state <= 7'd94;
wire _guard2681 = _guard2679 & _guard2680;
wire _guard2682 = ev00__0state >= 7'd94;
wire _guard2683 = ev00__0state <= 7'd94;
wire _guard2684 = _guard2682 & _guard2683;
wire _guard2685 = ev00__0state >= 7'd94;
wire _guard2686 = ev00__0state <= 7'd94;
wire _guard2687 = _guard2685 & _guard2686;
wire _guard2688 = ev00__0state >= 7'd94;
wire _guard2689 = ev00__0state <= 7'd94;
wire _guard2690 = _guard2688 & _guard2689;
wire _guard2691 = ev00__0state >= 7'd94;
wire _guard2692 = ev00__0state <= 7'd94;
wire _guard2693 = _guard2691 & _guard2692;
wire _guard2694 = ev00__0state >= 7'd94;
wire _guard2695 = ev00__0state <= 7'd94;
wire _guard2696 = _guard2694 & _guard2695;
wire _guard2697 = ev00__0state >= 7'd94;
wire _guard2698 = ev00__0state <= 7'd94;
wire _guard2699 = _guard2697 & _guard2698;
wire _guard2700 = ev00__0state >= 7'd94;
wire _guard2701 = ev00__0state <= 7'd94;
wire _guard2702 = _guard2700 & _guard2701;
wire _guard2703 = ev00__0state >= 7'd94;
wire _guard2704 = ev00__0state <= 7'd94;
wire _guard2705 = _guard2703 & _guard2704;
wire _guard2706 = ev00__0state >= 7'd94;
wire _guard2707 = ev00__0state <= 7'd94;
wire _guard2708 = _guard2706 & _guard2707;
wire _guard2709 = ev00__0state >= 7'd94;
wire _guard2710 = ev00__0state <= 7'd94;
wire _guard2711 = _guard2709 & _guard2710;
wire _guard2712 = ev00__0state >= 7'd94;
wire _guard2713 = ev00__0state <= 7'd94;
wire _guard2714 = _guard2712 & _guard2713;
wire _guard2715 = ev00__0state >= 7'd94;
wire _guard2716 = ev00__0state <= 7'd94;
wire _guard2717 = _guard2715 & _guard2716;
wire _guard2718 = ev00__0state >= 7'd94;
wire _guard2719 = ev00__0state <= 7'd94;
wire _guard2720 = _guard2718 & _guard2719;
wire _guard2721 = ev00__0state >= 7'd94;
wire _guard2722 = ev00__0state <= 7'd94;
wire _guard2723 = _guard2721 & _guard2722;
wire _guard2724 = ev00__0state >= 7'd94;
wire _guard2725 = ev00__0state <= 7'd94;
wire _guard2726 = _guard2724 & _guard2725;
wire _guard2727 = ev00__0state >= 7'd94;
wire _guard2728 = ev00__0state <= 7'd94;
wire _guard2729 = _guard2727 & _guard2728;
wire _guard2730 = ev00__0state >= 7'd94;
wire _guard2731 = ev00__0state <= 7'd94;
wire _guard2732 = _guard2730 & _guard2731;
wire _guard2733 = ev00__0state >= 7'd94;
wire _guard2734 = ev00__0state <= 7'd94;
wire _guard2735 = _guard2733 & _guard2734;
wire _guard2736 = ev00__0state >= 7'd94;
wire _guard2737 = ev00__0state <= 7'd94;
wire _guard2738 = _guard2736 & _guard2737;
wire _guard2739 = ev00__0state >= 7'd94;
wire _guard2740 = ev00__0state <= 7'd94;
wire _guard2741 = _guard2739 & _guard2740;
wire _guard2742 = ev00__0state >= 7'd94;
wire _guard2743 = ev00__0state <= 7'd94;
wire _guard2744 = _guard2742 & _guard2743;
wire _guard2745 = ev00__0state >= 7'd94;
wire _guard2746 = ev00__0state <= 7'd94;
wire _guard2747 = _guard2745 & _guard2746;
wire _guard2748 = ev00__0state >= 7'd94;
wire _guard2749 = ev00__0state <= 7'd94;
wire _guard2750 = _guard2748 & _guard2749;
wire _guard2751 = ev00__1_0;
wire _guard2752 = ev00__1state >= 7'd1;
wire _guard2753 = ev00__1state <= 7'd0;
wire _guard2754 = _guard2752 & _guard2753;
wire _guard2755 = _guard2751 | _guard2754;
wire _guard2756 = ev00__0state >= 7'd32;
wire _guard2757 = ev00__0state <= 7'd32;
wire _guard2758 = _guard2756 & _guard2757;
wire _guard2759 = ev00__0state >= 7'd64;
wire _guard2760 = ev00__0state <= 7'd64;
wire _guard2761 = _guard2759 & _guard2760;
wire _guard2762 = ev00__0state >= 7'd96;
wire _guard2763 = ev00__0state <= 7'd96;
wire _guard2764 = _guard2762 & _guard2763;
wire _guard2765 = ev00__0state >= 7'd31;
wire _guard2766 = ev00__0state <= 7'd31;
wire _guard2767 = _guard2765 & _guard2766;
wire _guard2768 = ev00__0state >= 7'd31;
wire _guard2769 = ev00__0state <= 7'd31;
wire _guard2770 = _guard2768 & _guard2769;
wire _guard2771 = ev00__0state >= 7'd31;
wire _guard2772 = ev00__0state <= 7'd31;
wire _guard2773 = _guard2771 & _guard2772;
wire _guard2774 = ev00__0state >= 7'd31;
wire _guard2775 = ev00__0state <= 7'd31;
wire _guard2776 = _guard2774 & _guard2775;
wire _guard2777 = ev00__0state >= 7'd31;
wire _guard2778 = ev00__0state <= 7'd31;
wire _guard2779 = _guard2777 & _guard2778;
wire _guard2780 = ev00__0state >= 7'd31;
wire _guard2781 = ev00__0state <= 7'd31;
wire _guard2782 = _guard2780 & _guard2781;
wire _guard2783 = ev00__0state >= 7'd31;
wire _guard2784 = ev00__0state <= 7'd31;
wire _guard2785 = _guard2783 & _guard2784;
wire _guard2786 = ev00__0state >= 7'd31;
wire _guard2787 = ev00__0state <= 7'd31;
wire _guard2788 = _guard2786 & _guard2787;
wire _guard2789 = ev00__0state >= 7'd31;
wire _guard2790 = ev00__0state <= 7'd31;
wire _guard2791 = _guard2789 & _guard2790;
wire _guard2792 = ev00__0state >= 7'd31;
wire _guard2793 = ev00__0state <= 7'd31;
wire _guard2794 = _guard2792 & _guard2793;
wire _guard2795 = ev00__0state >= 7'd31;
wire _guard2796 = ev00__0state <= 7'd31;
wire _guard2797 = _guard2795 & _guard2796;
wire _guard2798 = ev00__0state >= 7'd31;
wire _guard2799 = ev00__0state <= 7'd31;
wire _guard2800 = _guard2798 & _guard2799;
wire _guard2801 = ev00__0state >= 7'd31;
wire _guard2802 = ev00__0state <= 7'd31;
wire _guard2803 = _guard2801 & _guard2802;
wire _guard2804 = ev00__0state >= 7'd31;
wire _guard2805 = ev00__0state <= 7'd31;
wire _guard2806 = _guard2804 & _guard2805;
wire _guard2807 = ev00__0state >= 7'd31;
wire _guard2808 = ev00__0state <= 7'd31;
wire _guard2809 = _guard2807 & _guard2808;
wire _guard2810 = ev00__0state >= 7'd31;
wire _guard2811 = ev00__0state <= 7'd31;
wire _guard2812 = _guard2810 & _guard2811;
wire _guard2813 = ev00__0state >= 7'd31;
wire _guard2814 = ev00__0state <= 7'd31;
wire _guard2815 = _guard2813 & _guard2814;
wire _guard2816 = ev00__0state >= 7'd31;
wire _guard2817 = ev00__0state <= 7'd31;
wire _guard2818 = _guard2816 & _guard2817;
wire _guard2819 = ev00__0state >= 7'd31;
wire _guard2820 = ev00__0state <= 7'd31;
wire _guard2821 = _guard2819 & _guard2820;
wire _guard2822 = ev00__0state >= 7'd31;
wire _guard2823 = ev00__0state <= 7'd31;
wire _guard2824 = _guard2822 & _guard2823;
wire _guard2825 = ev00__0state >= 7'd31;
wire _guard2826 = ev00__0state <= 7'd31;
wire _guard2827 = _guard2825 & _guard2826;
wire _guard2828 = ev00__0state >= 7'd31;
wire _guard2829 = ev00__0state <= 7'd31;
wire _guard2830 = _guard2828 & _guard2829;
wire _guard2831 = ev00__0state >= 7'd31;
wire _guard2832 = ev00__0state <= 7'd31;
wire _guard2833 = _guard2831 & _guard2832;
wire _guard2834 = ev00__0state >= 7'd31;
wire _guard2835 = ev00__0state <= 7'd31;
wire _guard2836 = _guard2834 & _guard2835;
wire _guard2837 = ev00__0state >= 7'd31;
wire _guard2838 = ev00__0state <= 7'd31;
wire _guard2839 = _guard2837 & _guard2838;
wire _guard2840 = ev00__0state >= 7'd31;
wire _guard2841 = ev00__0state <= 7'd31;
wire _guard2842 = _guard2840 & _guard2841;
wire _guard2843 = ev00__0state >= 7'd31;
wire _guard2844 = ev00__0state <= 7'd31;
wire _guard2845 = _guard2843 & _guard2844;
wire _guard2846 = ev00__0state >= 7'd31;
wire _guard2847 = ev00__0state <= 7'd31;
wire _guard2848 = _guard2846 & _guard2847;
wire _guard2849 = ev00__0state >= 7'd31;
wire _guard2850 = ev00__0state <= 7'd31;
wire _guard2851 = _guard2849 & _guard2850;
wire _guard2852 = ev00__0state >= 7'd31;
wire _guard2853 = ev00__0state <= 7'd31;
wire _guard2854 = _guard2852 & _guard2853;
wire _guard2855 = ev00__0state >= 7'd31;
wire _guard2856 = ev00__0state <= 7'd31;
wire _guard2857 = _guard2855 & _guard2856;
wire _guard2858 = ev00__0state >= 7'd31;
wire _guard2859 = ev00__0state <= 7'd31;
wire _guard2860 = _guard2858 & _guard2859;
wire _guard2861 = ev00__0state >= 7'd127;
wire _guard2862 = ev00__0state <= 7'd127;
wire _guard2863 = _guard2861 & _guard2862;
wire _guard2864 = ev00__0state >= 7'd63;
wire _guard2865 = ev00__0state <= 7'd63;
wire _guard2866 = _guard2864 & _guard2865;
wire _guard2867 = ev00__0state >= 7'd95;
wire _guard2868 = ev00__0state <= 7'd95;
wire _guard2869 = _guard2867 & _guard2868;
wire _guard2870 = ev00__0state >= 7'd31;
wire _guard2871 = ev00__0state <= 7'd31;
wire _guard2872 = _guard2870 & _guard2871;
wire _guard2873 = ev00__0_0;
wire _guard2874 = ev00__0state >= 7'd1;
wire _guard2875 = ev00__0state <= 7'd0;
wire _guard2876 = _guard2874 & _guard2875;
wire _guard2877 = _guard2873 | _guard2876;
wire _guard2878 = ev00__0_0;
wire _guard2879 = ev00__0state >= 7'd1;
wire _guard2880 = ev00__0state <= 7'd0;
wire _guard2881 = _guard2879 & _guard2880;
wire _guard2882 = _guard2878 | _guard2881;
wire _guard2883 = ev00__0_0;
wire _guard2884 = ev00__0state >= 7'd1;
wire _guard2885 = ev00__0state <= 7'd0;
wire _guard2886 = _guard2884 & _guard2885;
wire _guard2887 = _guard2883 | _guard2886;
wire _guard2888 = ev00__0_0;
wire _guard2889 = ev00__0state >= 7'd1;
wire _guard2890 = ev00__0state <= 7'd0;
wire _guard2891 = _guard2889 & _guard2890;
wire _guard2892 = _guard2888 | _guard2891;
wire _guard2893 = ev00__0_0;
wire _guard2894 = ev00__0state >= 7'd1;
wire _guard2895 = ev00__0state <= 7'd0;
wire _guard2896 = _guard2894 & _guard2895;
wire _guard2897 = _guard2893 | _guard2896;
wire _guard2898 = ev00__0_0;
wire _guard2899 = ev00__0state >= 7'd1;
wire _guard2900 = ev00__0state <= 7'd0;
wire _guard2901 = _guard2899 & _guard2900;
wire _guard2902 = _guard2898 | _guard2901;
wire _guard2903 = ev00__0_0;
wire _guard2904 = ev00__0state >= 7'd1;
wire _guard2905 = ev00__0state <= 7'd0;
wire _guard2906 = _guard2904 & _guard2905;
wire _guard2907 = _guard2903 | _guard2906;
wire _guard2908 = ev00__0_0;
wire _guard2909 = ev00__0state >= 7'd1;
wire _guard2910 = ev00__0state <= 7'd0;
wire _guard2911 = _guard2909 & _guard2910;
wire _guard2912 = _guard2908 | _guard2911;
wire _guard2913 = ev00__0_0;
wire _guard2914 = ev00__0state >= 7'd1;
wire _guard2915 = ev00__0state <= 7'd0;
wire _guard2916 = _guard2914 & _guard2915;
wire _guard2917 = _guard2913 | _guard2916;
wire _guard2918 = ev00__0_0;
wire _guard2919 = ev00__0state >= 7'd1;
wire _guard2920 = ev00__0state <= 7'd0;
wire _guard2921 = _guard2919 & _guard2920;
wire _guard2922 = _guard2918 | _guard2921;
wire _guard2923 = ev00__0_0;
wire _guard2924 = ev00__0state >= 7'd1;
wire _guard2925 = ev00__0state <= 7'd0;
wire _guard2926 = _guard2924 & _guard2925;
wire _guard2927 = _guard2923 | _guard2926;
wire _guard2928 = ev00__0_0;
wire _guard2929 = ev00__0state >= 7'd1;
wire _guard2930 = ev00__0state <= 7'd0;
wire _guard2931 = _guard2929 & _guard2930;
wire _guard2932 = _guard2928 | _guard2931;
wire _guard2933 = ev00__0_0;
wire _guard2934 = ev00__0state >= 7'd1;
wire _guard2935 = ev00__0state <= 7'd0;
wire _guard2936 = _guard2934 & _guard2935;
wire _guard2937 = _guard2933 | _guard2936;
wire _guard2938 = ev00__0_0;
wire _guard2939 = ev00__0state >= 7'd1;
wire _guard2940 = ev00__0state <= 7'd0;
wire _guard2941 = _guard2939 & _guard2940;
wire _guard2942 = _guard2938 | _guard2941;
wire _guard2943 = ev00__0_0;
wire _guard2944 = ev00__0state >= 7'd1;
wire _guard2945 = ev00__0state <= 7'd0;
wire _guard2946 = _guard2944 & _guard2945;
wire _guard2947 = _guard2943 | _guard2946;
wire _guard2948 = ev00__0_0;
wire _guard2949 = ev00__0state >= 7'd1;
wire _guard2950 = ev00__0state <= 7'd0;
wire _guard2951 = _guard2949 & _guard2950;
wire _guard2952 = _guard2948 | _guard2951;
wire _guard2953 = ev00__0_0;
wire _guard2954 = ev00__0state >= 7'd1;
wire _guard2955 = ev00__0state <= 7'd0;
wire _guard2956 = _guard2954 & _guard2955;
wire _guard2957 = _guard2953 | _guard2956;
wire _guard2958 = ev00__0_0;
wire _guard2959 = ev00__0state >= 7'd1;
wire _guard2960 = ev00__0state <= 7'd0;
wire _guard2961 = _guard2959 & _guard2960;
wire _guard2962 = _guard2958 | _guard2961;
wire _guard2963 = ev00__0_0;
wire _guard2964 = ev00__0state >= 7'd1;
wire _guard2965 = ev00__0state <= 7'd0;
wire _guard2966 = _guard2964 & _guard2965;
wire _guard2967 = _guard2963 | _guard2966;
wire _guard2968 = ev00__0_0;
wire _guard2969 = ev00__0state >= 7'd1;
wire _guard2970 = ev00__0state <= 7'd0;
wire _guard2971 = _guard2969 & _guard2970;
wire _guard2972 = _guard2968 | _guard2971;
wire _guard2973 = ev00__0_0;
wire _guard2974 = ev00__0state >= 7'd1;
wire _guard2975 = ev00__0state <= 7'd0;
wire _guard2976 = _guard2974 & _guard2975;
wire _guard2977 = _guard2973 | _guard2976;
wire _guard2978 = ev00__0_0;
wire _guard2979 = ev00__0state >= 7'd1;
wire _guard2980 = ev00__0state <= 7'd0;
wire _guard2981 = _guard2979 & _guard2980;
wire _guard2982 = _guard2978 | _guard2981;
wire _guard2983 = ev00__0_0;
wire _guard2984 = ev00__0state >= 7'd1;
wire _guard2985 = ev00__0state <= 7'd0;
wire _guard2986 = _guard2984 & _guard2985;
wire _guard2987 = _guard2983 | _guard2986;
wire _guard2988 = ev00__0_0;
wire _guard2989 = ev00__0state >= 7'd1;
wire _guard2990 = ev00__0state <= 7'd0;
wire _guard2991 = _guard2989 & _guard2990;
wire _guard2992 = _guard2988 | _guard2991;
wire _guard2993 = ev00__0_0;
wire _guard2994 = ev00__0state >= 7'd1;
wire _guard2995 = ev00__0state <= 7'd0;
wire _guard2996 = _guard2994 & _guard2995;
wire _guard2997 = _guard2993 | _guard2996;
wire _guard2998 = ev00__0_0;
wire _guard2999 = ev00__0state >= 7'd1;
wire _guard3000 = ev00__0state <= 7'd0;
wire _guard3001 = _guard2999 & _guard3000;
wire _guard3002 = _guard2998 | _guard3001;
wire _guard3003 = ev00__0_0;
wire _guard3004 = ev00__0state >= 7'd1;
wire _guard3005 = ev00__0state <= 7'd0;
wire _guard3006 = _guard3004 & _guard3005;
wire _guard3007 = _guard3003 | _guard3006;
wire _guard3008 = ev00__0_0;
wire _guard3009 = ev00__0state >= 7'd1;
wire _guard3010 = ev00__0state <= 7'd0;
wire _guard3011 = _guard3009 & _guard3010;
wire _guard3012 = _guard3008 | _guard3011;
wire _guard3013 = ev00__0_0;
wire _guard3014 = ev00__0state >= 7'd1;
wire _guard3015 = ev00__0state <= 7'd0;
wire _guard3016 = _guard3014 & _guard3015;
wire _guard3017 = _guard3013 | _guard3016;
wire _guard3018 = ev00__0_0;
wire _guard3019 = ev00__0state >= 7'd1;
wire _guard3020 = ev00__0state <= 7'd0;
wire _guard3021 = _guard3019 & _guard3020;
wire _guard3022 = _guard3018 | _guard3021;
wire _guard3023 = ev00__0_0;
wire _guard3024 = ev00__0state >= 7'd1;
wire _guard3025 = ev00__0state <= 7'd0;
wire _guard3026 = _guard3024 & _guard3025;
wire _guard3027 = _guard3023 | _guard3026;
wire _guard3028 = ev00__0_0;
wire _guard3029 = ev00__0state >= 7'd1;
wire _guard3030 = ev00__0state <= 7'd0;
wire _guard3031 = _guard3029 & _guard3030;
wire _guard3032 = _guard3028 | _guard3031;
wire _guard3033 = ev00__0_0;
wire _guard3034 = ev00__0state >= 7'd1;
wire _guard3035 = ev00__0state <= 7'd0;
wire _guard3036 = _guard3034 & _guard3035;
wire _guard3037 = _guard3033 | _guard3036;
wire _guard3038 = ev00__0state >= 7'd31;
wire _guard3039 = ev00__0state <= 7'd31;
wire _guard3040 = _guard3038 & _guard3039;
assign p162 =
  _guard5 ? inst33_p27 :
  32'd0;
assign p167 =
  _guard10 ? inst33_p32 :
  32'd0;
assign p141 =
  _guard15 ? inst33_p6 :
  32'd0;
assign p143 =
  _guard20 ? inst33_p8 :
  32'd0;
assign p148 =
  _guard25 ? inst33_p13 :
  32'd0;
assign p161 =
  _guard30 ? inst33_p26 :
  32'd0;
assign p156 =
  _guard35 ? inst33_p21 :
  32'd0;
assign p157 =
  _guard40 ? inst33_p22 :
  32'd0;
assign p142 =
  _guard45 ? inst33_p7 :
  32'd0;
assign p168 =
  _guard50 ? inst33_p33 :
  32'd0;
assign p147 =
  _guard55 ? inst33_p12 :
  32'd0;
assign p169 =
  _guard60 ? inst33_p34 :
  32'd0;
assign p171 =
  _guard65 ? inst33_p36 :
  32'd0;
assign p155 =
  _guard70 ? inst33_p20 :
  32'd0;
assign p158 =
  _guard75 ? inst33_p23 :
  32'd0;
assign p170 =
  _guard80 ? inst33_p35 :
  32'd0;
assign p144 =
  _guard85 ? inst33_p9 :
  32'd0;
assign p163 =
  _guard90 ? inst33_p28 :
  32'd0;
assign p140 =
  _guard95 ? inst33_p5 :
  32'd0;
assign p149 =
  _guard100 ? inst33_p14 :
  32'd0;
assign p153 =
  _guard105 ? inst33_p18 :
  32'd0;
assign p165 =
  _guard110 ? inst33_p30 :
  32'd0;
assign p166 =
  _guard115 ? inst33_p31 :
  32'd0;
assign p145 =
  _guard120 ? inst33_p10 :
  32'd0;
assign p151 =
  _guard125 ? inst33_p16 :
  32'd0;
assign p154 =
  _guard130 ? inst33_p19 :
  32'd0;
assign p164 =
  _guard135 ? inst33_p29 :
  32'd0;
assign p150 =
  _guard140 ? inst33_p15 :
  32'd0;
assign p159 =
  _guard145 ? inst33_p24 :
  32'd0;
assign p160 =
  _guard150 ? inst33_p25 :
  32'd0;
assign p146 =
  _guard155 ? inst33_p11 :
  32'd0;
assign p152 =
  _guard160 ? inst33_p17 :
  32'd0;
assign inst5_p12 = inst2_p27;
assign inst5_p16 = inst2_p31;
assign inst5_p4 = inst2_p19;
assign inst5_p6 = inst2_p21;
assign inst5_p9 = inst2_p24;
assign inst5_p15 = inst2_p30;
assign inst5_p17 = inst2_p32;
assign inst5_clk = clk;
assign inst5_p11 = inst2_p26;
assign inst5_p5 = inst2_p20;
assign inst5_p8 = inst2_p23;
assign inst5_p10 = inst2_p25;
assign inst5_p2 = inst2_p17;
assign inst5_p3 = inst2_p18;
assign inst5_reset = reset;
assign inst5_p13 = inst2_p28;
assign inst5_p7 = inst2_p22;
assign inst5_p14 = inst2_p29;
assign inst21_p4 = inst9_out;
assign inst21_clk = clk;
assign inst21_reset = reset;
assign inst15_p19 = inst27_p19;
assign inst15_p28 = inst27_p28;
assign inst15_p29 = inst27_p29;
assign inst15_p12 = inst27_p12;
assign inst15_p16 = inst27_p16;
assign inst15_p6 = inst27_p6;
assign inst15_p9 = inst27_p9;
assign inst15_p15 = inst27_p15;
assign inst15_p17 = inst27_p17;
assign inst15_p20 = inst27_p20;
assign inst15_p21 = inst27_p21;
assign inst15_p23 = inst27_p23;
assign inst15_clk = clk;
assign inst15_p11 = inst27_p11;
assign inst15_p25 = inst27_p25;
assign inst15_p36 = inst27_p36;
assign inst15_p5 = inst27_p5;
assign inst15_p8 = inst27_p8;
assign inst15_p10 = inst27_p10;
assign inst15_reset = reset;
assign inst15_p13 = inst27_p13;
assign inst15_p18 = inst27_p18;
assign inst15_p30 = inst27_p30;
assign inst15_p7 = inst27_p7;
assign inst15_p24 = inst27_p24;
assign inst15_p32 = inst27_p32;
assign inst15_p14 = inst27_p14;
assign inst15_p26 = inst27_p26;
assign inst15_p31 = inst27_p31;
assign inst15_p27 = inst27_p27;
assign inst15_p33 = inst27_p33;
assign inst15_p22 = inst27_p22;
assign inst15_p34 = inst27_p34;
assign inst15_p35 = inst27_p35;
assign inst16_p19 = inst0_p105;
assign inst16_p28 = inst0_p114;
assign inst16_p29 = inst0_p115;
assign inst16_p12 = inst0_p98;
assign inst16_p16 = inst0_p102;
assign inst16_p6 = inst0_p92;
assign inst16_p9 = inst0_p95;
assign inst16_p15 = inst0_p101;
assign inst16_p17 = inst0_p103;
assign inst16_p20 = inst0_p106;
assign inst16_p21 = inst0_p107;
assign inst16_p23 = inst0_p109;
assign inst16_clk = clk;
assign inst16_p11 = inst0_p97;
assign inst16_p25 = inst0_p111;
assign inst16_p36 = inst0_p122;
assign inst16_p5 = inst0_p91;
assign inst16_p8 = inst0_p94;
assign inst16_p10 = inst0_p96;
assign inst16_reset = reset;
assign inst16_p13 = inst0_p99;
assign inst16_p18 = inst0_p104;
assign inst16_p30 = inst0_p116;
assign inst16_p7 = inst0_p93;
assign inst16_p24 = inst0_p110;
assign inst16_p32 = inst0_p118;
assign inst16_p14 = inst0_p100;
assign inst16_p26 = inst0_p112;
assign inst16_p31 = inst0_p117;
assign inst16_p27 = inst0_p113;
assign inst16_p33 = inst0_p119;
assign inst16_p22 = inst0_p108;
assign inst16_p34 = inst0_p120;
assign inst16_p35 = inst0_p121;
assign inst8_p12 = inst2_p27;
assign inst8_p16 = inst2_p31;
assign inst8_p4 = inst2_p19;
assign inst8_p6 = inst2_p21;
assign inst8_p9 = inst2_p24;
assign inst8_p15 = inst2_p30;
assign inst8_p17 = inst2_p32;
assign inst8_clk = clk;
assign inst8_p11 = inst2_p26;
assign inst8_p5 = inst2_p20;
assign inst8_p8 = inst2_p23;
assign inst8_p10 = inst2_p25;
assign inst8_p2 = inst2_p17;
assign inst8_p3 = inst2_p18;
assign inst8_reset = reset;
assign inst8_p13 = inst2_p28;
assign inst8_p7 = inst2_p22;
assign inst8_p14 = inst2_p29;
assign inst12_p19 = inst0_p105;
assign inst12_p28 = inst0_p114;
assign inst12_p29 = inst0_p115;
assign inst12_p12 = inst0_p98;
assign inst12_p16 = inst0_p102;
assign inst12_p6 = inst0_p92;
assign inst12_p9 = inst0_p95;
assign inst12_p15 = inst0_p101;
assign inst12_p17 = inst0_p103;
assign inst12_p20 = inst0_p106;
assign inst12_p21 = inst0_p107;
assign inst12_p23 = inst0_p109;
assign inst12_clk = clk;
assign inst12_p11 = inst0_p97;
assign inst12_p25 = inst0_p111;
assign inst12_p36 = inst0_p122;
assign inst12_p5 = inst0_p91;
assign inst12_p8 = inst0_p94;
assign inst12_p10 = inst0_p96;
assign inst12_reset = reset;
assign inst12_p13 = inst0_p99;
assign inst12_p18 = inst0_p104;
assign inst12_p30 = inst0_p116;
assign inst12_p7 = inst0_p93;
assign inst12_p24 = inst0_p110;
assign inst12_p32 = inst0_p118;
assign inst12_p14 = inst0_p100;
assign inst12_p26 = inst0_p112;
assign inst12_p31 = inst0_p117;
assign inst12_p27 = inst0_p113;
assign inst12_p33 = inst0_p119;
assign inst12_p22 = inst0_p108;
assign inst12_p34 = inst0_p120;
assign inst12_p35 = inst0_p121;
assign inst31_p4 = inst4_out;
assign inst31_clk = clk;
assign inst31_reset = reset;
assign inst32_p19 = inst1_p48;
assign inst32_p28 = inst1_p57;
assign inst32_p29 = inst1_p58;
assign inst32_p12 = inst1_p41;
assign inst32_p16 = inst1_p45;
assign inst32_p6 = inst1_p35;
assign inst32_p9 = inst1_p38;
assign inst32_p15 = inst1_p44;
assign inst32_p17 = inst1_p46;
assign inst32_p20 = inst1_p49;
assign inst32_p21 = inst1_p50;
assign inst32_p23 = inst1_p52;
assign inst32_clk = clk;
assign inst32_p11 = inst1_p40;
assign inst32_p25 = inst1_p54;
assign inst32_p36 = inst1_p65;
assign inst32_p5 = inst1_p34;
assign inst32_p8 = inst1_p37;
assign inst32_p10 = inst1_p39;
assign inst32_reset = reset;
assign inst32_p13 = inst1_p42;
assign inst32_p18 = inst1_p47;
assign inst32_p30 = inst1_p59;
assign inst32_p7 = inst1_p36;
assign inst32_p24 = inst1_p53;
assign inst32_p32 = inst1_p61;
assign inst32_p14 = inst1_p43;
assign inst32_p26 = inst1_p55;
assign inst32_p31 = inst1_p60;
assign inst32_p27 = inst1_p56;
assign inst32_p33 = inst1_p62;
assign inst32_p22 = inst1_p51;
assign inst32_p34 = inst1_p63;
assign inst32_p35 = inst1_p64;
assign inst3_p19 = p125;
assign inst3_p28 = p134;
assign inst3_p29 = p135;
assign inst3_p12 = p118;
assign inst3_p16 = p122;
assign inst3_p4 = p110;
assign inst3_p6 = p112;
assign inst3_p9 = p115;
assign inst3_p15 = p121;
assign inst3_p17 = p123;
assign inst3_p20 = p126;
assign inst3_p21 = p127;
assign inst3_p23 = p129;
assign inst3_clk = clk;
assign inst3_p11 = p117;
assign inst3_p25 = p131;
assign inst3_p5 = p111;
assign inst3_p8 = p114;
assign inst3_p10 = p116;
assign inst3_p2 = p108;
assign inst3_p3 = p109;
assign inst3_reset = reset;
assign inst3_p13 = p119;
assign inst3_p18 = p124;
assign inst3_p30 = p136;
assign inst3_p7 = p113;
assign inst3_p24 = p130;
assign inst3_p32 = p138;
assign inst3_p14 = p120;
assign inst3_p26 = p132;
assign inst3_p31 = p137;
assign inst3_p27 = p133;
assign inst3_p33 = p139;
assign inst3_p22 = p128;
assign inst25_p4 = inst9_out;
assign inst25_clk = clk;
assign inst25_reset = reset;
assign inst29_p4 = inst4_out;
assign inst29_clk = clk;
assign inst29_reset = reset;
assign inst28_p19 = inst1_p48;
assign inst28_p28 = inst1_p57;
assign inst28_p29 = inst1_p58;
assign inst28_p12 = inst1_p41;
assign inst28_p16 = inst1_p45;
assign inst28_p6 = inst1_p35;
assign inst28_p9 = inst1_p38;
assign inst28_p15 = inst1_p44;
assign inst28_p17 = inst1_p46;
assign inst28_p20 = inst1_p49;
assign inst28_p21 = inst1_p50;
assign inst28_p23 = inst1_p52;
assign inst28_clk = clk;
assign inst28_p11 = inst1_p40;
assign inst28_p25 = inst1_p54;
assign inst28_p36 = inst1_p65;
assign inst28_p5 = inst1_p34;
assign inst28_p8 = inst1_p37;
assign inst28_p10 = inst1_p39;
assign inst28_reset = reset;
assign inst28_p13 = inst1_p42;
assign inst28_p18 = inst1_p47;
assign inst28_p30 = inst1_p59;
assign inst28_p7 = inst1_p36;
assign inst28_p24 = inst1_p53;
assign inst28_p32 = inst1_p61;
assign inst28_p14 = inst1_p43;
assign inst28_p26 = inst1_p55;
assign inst28_p31 = inst1_p60;
assign inst28_p27 = inst1_p56;
assign inst28_p33 = inst1_p62;
assign inst28_p22 = inst1_p51;
assign inst28_p34 = inst1_p63;
assign inst28_p35 = inst1_p64;
assign inst9_write_en = _guard1005;
assign inst9_clk = clk;
assign inst9_reset = reset;
assign inst9_in =
  _guard1008 ? inst15_p37 :
  _guard1011 ? inst16_p37 :
  _guard1014 ? inst12_p37 :
  _guard1017 ? inst24_p37 :
  _guard1020 ? inst23_p37 :
  _guard1023 ? inst19_p37 :
  _guard1026 ? inst20_p37 :
  _guard1031 ? inst11_p37 :
  'x;
assign inst17_p4 = inst9_out;
assign inst17_clk = clk;
assign inst17_reset = reset;
assign inst1_p19 =
  _guard1037 ? inst21_p22 :
  _guard1040 ? inst25_p22 :
  _guard1043 ? inst17_p22 :
  _guard1046 ? inst13_p22 :
  'x;
assign inst1_p28 =
  _guard1049 ? inst21_p31 :
  _guard1052 ? inst25_p31 :
  _guard1055 ? inst17_p31 :
  _guard1058 ? inst13_p31 :
  'x;
assign inst1_p29 =
  _guard1061 ? inst21_p32 :
  _guard1064 ? inst25_p32 :
  _guard1067 ? inst17_p32 :
  _guard1070 ? inst13_p32 :
  'x;
assign inst1_p12 =
  _guard1073 ? inst21_p15 :
  _guard1076 ? inst25_p15 :
  _guard1079 ? inst17_p15 :
  _guard1082 ? inst13_p15 :
  'x;
assign inst1_p16 =
  _guard1085 ? inst21_p19 :
  _guard1088 ? inst25_p19 :
  _guard1091 ? inst17_p19 :
  _guard1094 ? inst13_p19 :
  'x;
assign inst1_p4 =
  _guard1097 ? inst21_p7 :
  _guard1100 ? inst25_p7 :
  _guard1103 ? inst17_p7 :
  _guard1106 ? inst13_p7 :
  'x;
assign inst1_p6 =
  _guard1109 ? inst21_p9 :
  _guard1112 ? inst25_p9 :
  _guard1115 ? inst17_p9 :
  _guard1118 ? inst13_p9 :
  'x;
assign inst1_p9 =
  _guard1121 ? inst21_p12 :
  _guard1124 ? inst25_p12 :
  _guard1127 ? inst17_p12 :
  _guard1130 ? inst13_p12 :
  'x;
assign inst1_p15 =
  _guard1133 ? inst21_p18 :
  _guard1136 ? inst25_p18 :
  _guard1139 ? inst17_p18 :
  _guard1142 ? inst13_p18 :
  'x;
assign inst1_p17 =
  _guard1145 ? inst21_p20 :
  _guard1148 ? inst25_p20 :
  _guard1151 ? inst17_p20 :
  _guard1154 ? inst13_p20 :
  'x;
assign inst1_p20 =
  _guard1157 ? inst21_p23 :
  _guard1160 ? inst25_p23 :
  _guard1163 ? inst17_p23 :
  _guard1166 ? inst13_p23 :
  'x;
assign inst1_p21 =
  _guard1169 ? inst21_p24 :
  _guard1172 ? inst25_p24 :
  _guard1175 ? inst17_p24 :
  _guard1178 ? inst13_p24 :
  'x;
assign inst1_p23 =
  _guard1181 ? inst21_p26 :
  _guard1184 ? inst25_p26 :
  _guard1187 ? inst17_p26 :
  _guard1190 ? inst13_p26 :
  'x;
assign inst1_clk = clk;
assign inst1_p11 =
  _guard1193 ? inst21_p14 :
  _guard1196 ? inst25_p14 :
  _guard1199 ? inst17_p14 :
  _guard1202 ? inst13_p14 :
  'x;
assign inst1_p25 =
  _guard1205 ? inst21_p28 :
  _guard1208 ? inst25_p28 :
  _guard1211 ? inst17_p28 :
  _guard1214 ? inst13_p28 :
  'x;
assign inst1_p5 =
  _guard1217 ? inst21_p8 :
  _guard1220 ? inst25_p8 :
  _guard1223 ? inst17_p8 :
  _guard1226 ? inst13_p8 :
  'x;
assign inst1_p8 =
  _guard1229 ? inst21_p11 :
  _guard1232 ? inst25_p11 :
  _guard1235 ? inst17_p11 :
  _guard1238 ? inst13_p11 :
  'x;
assign inst1_p10 =
  _guard1241 ? inst21_p13 :
  _guard1244 ? inst25_p13 :
  _guard1247 ? inst17_p13 :
  _guard1250 ? inst13_p13 :
  'x;
assign inst1_p2 =
  _guard1253 ? inst21_p5 :
  _guard1256 ? inst25_p5 :
  _guard1259 ? inst17_p5 :
  _guard1262 ? inst13_p5 :
  'x;
assign inst1_p3 =
  _guard1265 ? inst21_p6 :
  _guard1268 ? inst25_p6 :
  _guard1271 ? inst17_p6 :
  _guard1274 ? inst13_p6 :
  'x;
assign inst1_reset = reset;
assign inst1_p13 =
  _guard1277 ? inst21_p16 :
  _guard1280 ? inst25_p16 :
  _guard1283 ? inst17_p16 :
  _guard1286 ? inst13_p16 :
  'x;
assign inst1_p18 =
  _guard1289 ? inst21_p21 :
  _guard1292 ? inst25_p21 :
  _guard1295 ? inst17_p21 :
  _guard1298 ? inst13_p21 :
  'x;
assign inst1_p30 =
  _guard1301 ? inst21_p33 :
  _guard1304 ? inst25_p33 :
  _guard1307 ? inst17_p33 :
  _guard1310 ? inst13_p33 :
  'x;
assign inst1_p7 =
  _guard1313 ? inst21_p10 :
  _guard1316 ? inst25_p10 :
  _guard1319 ? inst17_p10 :
  _guard1322 ? inst13_p10 :
  'x;
assign inst1_p24 =
  _guard1325 ? inst21_p27 :
  _guard1328 ? inst25_p27 :
  _guard1331 ? inst17_p27 :
  _guard1334 ? inst13_p27 :
  'x;
assign inst1_p32 =
  _guard1337 ? inst21_p35 :
  _guard1340 ? inst25_p35 :
  _guard1343 ? inst17_p35 :
  _guard1346 ? inst13_p35 :
  'x;
assign inst1_p14 =
  _guard1349 ? inst21_p17 :
  _guard1352 ? inst25_p17 :
  _guard1355 ? inst17_p17 :
  _guard1358 ? inst13_p17 :
  'x;
assign inst1_p26 =
  _guard1361 ? inst21_p29 :
  _guard1364 ? inst25_p29 :
  _guard1367 ? inst17_p29 :
  _guard1370 ? inst13_p29 :
  'x;
assign inst1_p31 =
  _guard1373 ? inst21_p34 :
  _guard1376 ? inst25_p34 :
  _guard1379 ? inst17_p34 :
  _guard1382 ? inst13_p34 :
  'x;
assign inst1_p27 =
  _guard1385 ? inst21_p30 :
  _guard1388 ? inst25_p30 :
  _guard1391 ? inst17_p30 :
  _guard1394 ? inst13_p30 :
  'x;
assign inst1_p33 =
  _guard1397 ? inst21_p36 :
  _guard1400 ? inst25_p36 :
  _guard1403 ? inst17_p36 :
  _guard1406 ? inst13_p36 :
  'x;
assign inst1_p22 =
  _guard1409 ? inst21_p25 :
  _guard1412 ? inst25_p25 :
  _guard1415 ? inst17_p25 :
  _guard1418 ? inst13_p25 :
  'x;
assign inst24_p19 = inst0_p105;
assign inst24_p28 = inst0_p114;
assign inst24_p29 = inst0_p115;
assign inst24_p12 = inst0_p98;
assign inst24_p16 = inst0_p102;
assign inst24_p6 = inst0_p92;
assign inst24_p9 = inst0_p95;
assign inst24_p15 = inst0_p101;
assign inst24_p17 = inst0_p103;
assign inst24_p20 = inst0_p106;
assign inst24_p21 = inst0_p107;
assign inst24_p23 = inst0_p109;
assign inst24_clk = clk;
assign inst24_p11 = inst0_p97;
assign inst24_p25 = inst0_p111;
assign inst24_p36 = inst0_p122;
assign inst24_p5 = inst0_p91;
assign inst24_p8 = inst0_p94;
assign inst24_p10 = inst0_p96;
assign inst24_reset = reset;
assign inst24_p13 = inst0_p99;
assign inst24_p18 = inst0_p104;
assign inst24_p30 = inst0_p116;
assign inst24_p7 = inst0_p93;
assign inst24_p24 = inst0_p110;
assign inst24_p32 = inst0_p118;
assign inst24_p14 = inst0_p100;
assign inst24_p26 = inst0_p112;
assign inst24_p31 = inst0_p117;
assign inst24_p27 = inst0_p113;
assign inst24_p33 = inst0_p119;
assign inst24_p22 = inst0_p108;
assign inst24_p34 = inst0_p120;
assign inst24_p35 = inst0_p121;
assign inst0_p47 =
  _guard1517 ? inst14_p9 :
  _guard1520 ? inst18_p9 :
  _guard1523 ? inst22_p9 :
  _guard1528 ? inst10_p9 :
  'x;
assign inst0_p70 =
  _guard1531 ? inst14_p32 :
  _guard1534 ? inst18_p32 :
  _guard1537 ? inst22_p32 :
  _guard1542 ? inst10_p32 :
  'x;
assign inst0_p80 =
  _guard1547 ? inst5_p23 :
  _guard1550 ? inst8_p23 :
  _guard1553 ? inst7_p23 :
  _guard1556 ? inst6_p23 :
  'x;
assign inst0_p65 =
  _guard1559 ? inst14_p27 :
  _guard1562 ? inst18_p27 :
  _guard1565 ? inst22_p27 :
  _guard1570 ? inst10_p27 :
  'x;
assign inst0_p74 =
  _guard1573 ? inst14_p36 :
  _guard1576 ? inst18_p36 :
  _guard1579 ? inst22_p36 :
  _guard1584 ? inst10_p36 :
  'x;
assign inst0_ev0 = _guard1601;
assign inst0_p52 =
  _guard1604 ? inst14_p14 :
  _guard1607 ? inst18_p14 :
  _guard1610 ? inst22_p14 :
  _guard1615 ? inst10_p14 :
  'x;
assign inst0_p59 =
  _guard1618 ? inst14_p21 :
  _guard1621 ? inst18_p21 :
  _guard1624 ? inst22_p21 :
  _guard1629 ? inst10_p21 :
  'x;
assign inst0_p56 =
  _guard1632 ? inst14_p18 :
  _guard1635 ? inst18_p18 :
  _guard1638 ? inst22_p18 :
  _guard1643 ? inst10_p18 :
  'x;
assign inst0_p68 =
  _guard1646 ? inst14_p30 :
  _guard1649 ? inst18_p30 :
  _guard1652 ? inst22_p30 :
  _guard1657 ? inst10_p30 :
  'x;
assign inst0_p79 =
  _guard1662 ? inst5_p22 :
  _guard1665 ? inst8_p22 :
  _guard1668 ? inst7_p22 :
  _guard1671 ? inst6_p22 :
  'x;
assign inst0_p60 =
  _guard1674 ? inst14_p22 :
  _guard1677 ? inst18_p22 :
  _guard1680 ? inst22_p22 :
  _guard1685 ? inst10_p22 :
  'x;
assign inst0_p64 =
  _guard1688 ? inst14_p26 :
  _guard1691 ? inst18_p26 :
  _guard1694 ? inst22_p26 :
  _guard1699 ? inst10_p26 :
  'x;
assign inst0_clk = clk;
assign inst0_p71 =
  _guard1702 ? inst14_p33 :
  _guard1705 ? inst18_p33 :
  _guard1708 ? inst22_p33 :
  _guard1713 ? inst10_p33 :
  'x;
assign inst0_p46 =
  _guard1716 ? inst14_p8 :
  _guard1719 ? inst18_p8 :
  _guard1722 ? inst22_p8 :
  _guard1727 ? inst10_p8 :
  'x;
assign inst0_p51 =
  _guard1730 ? inst14_p13 :
  _guard1733 ? inst18_p13 :
  _guard1736 ? inst22_p13 :
  _guard1741 ? inst10_p13 :
  'x;
assign inst0_p54 =
  _guard1744 ? inst14_p16 :
  _guard1747 ? inst18_p16 :
  _guard1750 ? inst22_p16 :
  _guard1755 ? inst10_p16 :
  'x;
assign inst0_p83 =
  _guard1760 ? inst5_p26 :
  _guard1763 ? inst8_p26 :
  _guard1766 ? inst7_p26 :
  _guard1769 ? inst6_p26 :
  'x;
assign inst0_p84 =
  _guard1774 ? inst5_p27 :
  _guard1777 ? inst8_p27 :
  _guard1780 ? inst7_p27 :
  _guard1783 ? inst6_p27 :
  'x;
assign inst0_p45 =
  _guard1786 ? inst14_p7 :
  _guard1789 ? inst18_p7 :
  _guard1792 ? inst22_p7 :
  _guard1797 ? inst10_p7 :
  'x;
assign inst0_p73 =
  _guard1800 ? inst14_p35 :
  _guard1803 ? inst18_p35 :
  _guard1806 ? inst22_p35 :
  _guard1811 ? inst10_p35 :
  'x;
assign inst0_p76 =
  _guard1816 ? inst5_p19 :
  _guard1819 ? inst8_p19 :
  _guard1822 ? inst7_p19 :
  _guard1825 ? inst6_p19 :
  'x;
assign inst0_p53 =
  _guard1828 ? inst14_p15 :
  _guard1831 ? inst18_p15 :
  _guard1834 ? inst22_p15 :
  _guard1839 ? inst10_p15 :
  'x;
assign inst0_p58 =
  _guard1842 ? inst14_p20 :
  _guard1845 ? inst18_p20 :
  _guard1848 ? inst22_p20 :
  _guard1853 ? inst10_p20 :
  'x;
assign inst0_p88 =
  _guard1858 ? inst5_p31 :
  _guard1861 ? inst8_p31 :
  _guard1864 ? inst7_p31 :
  _guard1867 ? inst6_p31 :
  'x;
assign inst0_p90 =
  _guard1872 ? inst5_p33 :
  _guard1875 ? inst8_p33 :
  _guard1878 ? inst7_p33 :
  _guard1881 ? inst6_p33 :
  'x;
assign inst0_reset = reset;
assign inst0_p50 =
  _guard1884 ? inst14_p12 :
  _guard1887 ? inst18_p12 :
  _guard1890 ? inst22_p12 :
  _guard1895 ? inst10_p12 :
  'x;
assign inst0_p75 =
  _guard1900 ? inst5_p18 :
  _guard1903 ? inst8_p18 :
  _guard1906 ? inst7_p18 :
  _guard1909 ? inst6_p18 :
  'x;
assign inst0_p43 =
  _guard1912 ? inst14_p5 :
  _guard1915 ? inst18_p5 :
  _guard1918 ? inst22_p5 :
  _guard1923 ? inst10_p5 :
  'x;
assign inst0_p72 =
  _guard1926 ? inst14_p34 :
  _guard1929 ? inst18_p34 :
  _guard1932 ? inst22_p34 :
  _guard1937 ? inst10_p34 :
  'x;
assign inst0_p77 =
  _guard1942 ? inst5_p20 :
  _guard1945 ? inst8_p20 :
  _guard1948 ? inst7_p20 :
  _guard1951 ? inst6_p20 :
  'x;
assign inst0_p63 =
  _guard1954 ? inst14_p25 :
  _guard1957 ? inst18_p25 :
  _guard1960 ? inst22_p25 :
  _guard1965 ? inst10_p25 :
  'x;
assign inst0_p69 =
  _guard1968 ? inst14_p31 :
  _guard1971 ? inst18_p31 :
  _guard1974 ? inst22_p31 :
  _guard1979 ? inst10_p31 :
  'x;
assign inst0_p87 =
  _guard1984 ? inst5_p30 :
  _guard1987 ? inst8_p30 :
  _guard1990 ? inst7_p30 :
  _guard1993 ? inst6_p30 :
  'x;
assign inst0_p89 =
  _guard1998 ? inst5_p32 :
  _guard2001 ? inst8_p32 :
  _guard2004 ? inst7_p32 :
  _guard2007 ? inst6_p32 :
  'x;
assign inst0_p48 =
  _guard2010 ? inst14_p10 :
  _guard2013 ? inst18_p10 :
  _guard2016 ? inst22_p10 :
  _guard2021 ? inst10_p10 :
  'x;
assign inst0_p49 =
  _guard2024 ? inst14_p11 :
  _guard2027 ? inst18_p11 :
  _guard2030 ? inst22_p11 :
  _guard2035 ? inst10_p11 :
  'x;
assign inst0_p61 =
  _guard2038 ? inst14_p23 :
  _guard2041 ? inst18_p23 :
  _guard2044 ? inst22_p23 :
  _guard2049 ? inst10_p23 :
  'x;
assign inst0_p81 =
  _guard2054 ? inst5_p24 :
  _guard2057 ? inst8_p24 :
  _guard2060 ? inst7_p24 :
  _guard2063 ? inst6_p24 :
  'x;
assign inst0_p62 =
  _guard2066 ? inst14_p24 :
  _guard2069 ? inst18_p24 :
  _guard2072 ? inst22_p24 :
  _guard2077 ? inst10_p24 :
  'x;
assign inst0_p66 =
  _guard2080 ? inst14_p28 :
  _guard2083 ? inst18_p28 :
  _guard2086 ? inst22_p28 :
  _guard2091 ? inst10_p28 :
  'x;
assign inst0_p85 =
  _guard2096 ? inst5_p28 :
  _guard2099 ? inst8_p28 :
  _guard2102 ? inst7_p28 :
  _guard2105 ? inst6_p28 :
  'x;
assign inst0_p57 =
  _guard2108 ? inst14_p19 :
  _guard2111 ? inst18_p19 :
  _guard2114 ? inst22_p19 :
  _guard2119 ? inst10_p19 :
  'x;
assign inst0_p78 =
  _guard2124 ? inst5_p21 :
  _guard2127 ? inst8_p21 :
  _guard2130 ? inst7_p21 :
  _guard2133 ? inst6_p21 :
  'x;
assign inst0_p82 =
  _guard2138 ? inst5_p25 :
  _guard2141 ? inst8_p25 :
  _guard2144 ? inst7_p25 :
  _guard2147 ? inst6_p25 :
  'x;
assign inst0_p44 =
  _guard2150 ? inst14_p6 :
  _guard2153 ? inst18_p6 :
  _guard2156 ? inst22_p6 :
  _guard2161 ? inst10_p6 :
  'x;
assign inst0_p55 =
  _guard2164 ? inst14_p17 :
  _guard2167 ? inst18_p17 :
  _guard2170 ? inst22_p17 :
  _guard2175 ? inst10_p17 :
  'x;
assign inst0_p67 =
  _guard2178 ? inst14_p29 :
  _guard2181 ? inst18_p29 :
  _guard2184 ? inst22_p29 :
  _guard2189 ? inst10_p29 :
  'x;
assign inst0_p86 =
  _guard2194 ? inst5_p29 :
  _guard2197 ? inst8_p29 :
  _guard2200 ? inst7_p29 :
  _guard2203 ? inst6_p29 :
  'x;
assign inst7_p12 = inst2_p27;
assign inst7_p16 = inst2_p31;
assign inst7_p4 = inst2_p19;
assign inst7_p6 = inst2_p21;
assign inst7_p9 = inst2_p24;
assign inst7_p15 = inst2_p30;
assign inst7_p17 = inst2_p32;
assign inst7_clk = clk;
assign inst7_p11 = inst2_p26;
assign inst7_p5 = inst2_p20;
assign inst7_p8 = inst2_p23;
assign inst7_p10 = inst2_p25;
assign inst7_p2 = inst2_p17;
assign inst7_p3 = inst2_p18;
assign inst7_reset = reset;
assign inst7_p13 = inst2_p28;
assign inst7_p7 = inst2_p22;
assign inst7_p14 = inst2_p29;
assign inst23_p19 = inst31_p19;
assign inst23_p28 = inst31_p28;
assign inst23_p29 = inst31_p29;
assign inst23_p12 = inst31_p12;
assign inst23_p16 = inst31_p16;
assign inst23_p6 = inst31_p6;
assign inst23_p9 = inst31_p9;
assign inst23_p15 = inst31_p15;
assign inst23_p17 = inst31_p17;
assign inst23_p20 = inst31_p20;
assign inst23_p21 = inst31_p21;
assign inst23_p23 = inst31_p23;
assign inst23_clk = clk;
assign inst23_p11 = inst31_p11;
assign inst23_p25 = inst31_p25;
assign inst23_p36 = inst31_p36;
assign inst23_p5 = inst31_p5;
assign inst23_p8 = inst31_p8;
assign inst23_p10 = inst31_p10;
assign inst23_reset = reset;
assign inst23_p13 = inst31_p13;
assign inst23_p18 = inst31_p18;
assign inst23_p30 = inst31_p30;
assign inst23_p7 = inst31_p7;
assign inst23_p24 = inst31_p24;
assign inst23_p32 = inst31_p32;
assign inst23_p14 = inst31_p14;
assign inst23_p26 = inst31_p26;
assign inst23_p31 = inst31_p31;
assign inst23_p27 = inst31_p27;
assign inst23_p33 = inst31_p33;
assign inst23_p22 = inst31_p22;
assign inst23_p34 = inst31_p34;
assign inst23_p35 = inst31_p35;
assign inst27_p4 = inst4_out;
assign inst27_clk = clk;
assign inst27_reset = reset;
assign inst30_p19 = inst1_p48;
assign inst30_p28 = inst1_p57;
assign inst30_p29 = inst1_p58;
assign inst30_p12 = inst1_p41;
assign inst30_p16 = inst1_p45;
assign inst30_p6 = inst1_p35;
assign inst30_p9 = inst1_p38;
assign inst30_p15 = inst1_p44;
assign inst30_p17 = inst1_p46;
assign inst30_p20 = inst1_p49;
assign inst30_p21 = inst1_p50;
assign inst30_p23 = inst1_p52;
assign inst30_clk = clk;
assign inst30_p11 = inst1_p40;
assign inst30_p25 = inst1_p54;
assign inst30_p36 = inst1_p65;
assign inst30_p5 = inst1_p34;
assign inst30_p8 = inst1_p37;
assign inst30_p10 = inst1_p39;
assign inst30_reset = reset;
assign inst30_p13 = inst1_p42;
assign inst30_p18 = inst1_p47;
assign inst30_p30 = inst1_p59;
assign inst30_p7 = inst1_p36;
assign inst30_p24 = inst1_p53;
assign inst30_p32 = inst1_p61;
assign inst30_p14 = inst1_p43;
assign inst30_p26 = inst1_p55;
assign inst30_p31 = inst1_p60;
assign inst30_p27 = inst1_p56;
assign inst30_p33 = inst1_p62;
assign inst30_p22 = inst1_p51;
assign inst30_p34 = inst1_p63;
assign inst30_p35 = inst1_p64;
assign inst19_p19 = inst29_p19;
assign inst19_p28 = inst29_p28;
assign inst19_p29 = inst29_p29;
assign inst19_p12 = inst29_p12;
assign inst19_p16 = inst29_p16;
assign inst19_p6 = inst29_p6;
assign inst19_p9 = inst29_p9;
assign inst19_p15 = inst29_p15;
assign inst19_p17 = inst29_p17;
assign inst19_p20 = inst29_p20;
assign inst19_p21 = inst29_p21;
assign inst19_p23 = inst29_p23;
assign inst19_clk = clk;
assign inst19_p11 = inst29_p11;
assign inst19_p25 = inst29_p25;
assign inst19_p36 = inst29_p36;
assign inst19_p5 = inst29_p5;
assign inst19_p8 = inst29_p8;
assign inst19_p10 = inst29_p10;
assign inst19_reset = reset;
assign inst19_p13 = inst29_p13;
assign inst19_p18 = inst29_p18;
assign inst19_p30 = inst29_p30;
assign inst19_p7 = inst29_p7;
assign inst19_p24 = inst29_p24;
assign inst19_p32 = inst29_p32;
assign inst19_p14 = inst29_p14;
assign inst19_p26 = inst29_p26;
assign inst19_p31 = inst29_p31;
assign inst19_p27 = inst29_p27;
assign inst19_p33 = inst29_p33;
assign inst19_p22 = inst29_p22;
assign inst19_p34 = inst29_p34;
assign inst19_p35 = inst29_p35;
assign ev00_clk = clk;
assign ev00_go = ev0;
assign ev00_reset = reset;
assign inst6_p12 = inst2_p27;
assign inst6_p16 = inst2_p31;
assign inst6_p4 = inst2_p19;
assign inst6_p6 = inst2_p21;
assign inst6_p9 = inst2_p24;
assign inst6_p15 = inst2_p30;
assign inst6_p17 = inst2_p32;
assign inst6_clk = clk;
assign inst6_p11 = inst2_p26;
assign inst6_p5 = inst2_p20;
assign inst6_p8 = inst2_p23;
assign inst6_p10 = inst2_p25;
assign inst6_p2 = inst2_p17;
assign inst6_p3 = inst2_p18;
assign inst6_reset = reset;
assign inst6_p13 = inst2_p28;
assign inst6_p7 = inst2_p22;
assign inst6_p14 = inst2_p29;
assign inst20_p19 = inst0_p105;
assign inst20_p28 = inst0_p114;
assign inst20_p29 = inst0_p115;
assign inst20_p12 = inst0_p98;
assign inst20_p16 = inst0_p102;
assign inst20_p6 = inst0_p92;
assign inst20_p9 = inst0_p95;
assign inst20_p15 = inst0_p101;
assign inst20_p17 = inst0_p103;
assign inst20_p20 = inst0_p106;
assign inst20_p21 = inst0_p107;
assign inst20_p23 = inst0_p109;
assign inst20_clk = clk;
assign inst20_p11 = inst0_p97;
assign inst20_p25 = inst0_p111;
assign inst20_p36 = inst0_p122;
assign inst20_p5 = inst0_p91;
assign inst20_p8 = inst0_p94;
assign inst20_p10 = inst0_p96;
assign inst20_reset = reset;
assign inst20_p13 = inst0_p99;
assign inst20_p18 = inst0_p104;
assign inst20_p30 = inst0_p116;
assign inst20_p7 = inst0_p93;
assign inst20_p24 = inst0_p110;
assign inst20_p32 = inst0_p118;
assign inst20_p14 = inst0_p100;
assign inst20_p26 = inst0_p112;
assign inst20_p31 = inst0_p117;
assign inst20_p27 = inst0_p113;
assign inst20_p33 = inst0_p119;
assign inst20_p22 = inst0_p108;
assign inst20_p34 = inst0_p120;
assign inst20_p35 = inst0_p121;
assign inst33_p4 = inst4_out;
assign inst33_clk = clk;
assign inst33_reset = reset;
assign inst14_p4 = inst9_out;
assign inst14_clk = clk;
assign inst14_reset = reset;
assign inst18_p4 = inst9_out;
assign inst18_clk = clk;
assign inst18_reset = reset;
assign inst22_p4 = inst9_out;
assign inst22_clk = clk;
assign inst22_reset = reset;
assign inst26_p19 = inst1_p48;
assign inst26_p28 = inst1_p57;
assign inst26_p29 = inst1_p58;
assign inst26_p12 = inst1_p41;
assign inst26_p16 = inst1_p45;
assign inst26_p6 = inst1_p35;
assign inst26_p9 = inst1_p38;
assign inst26_p15 = inst1_p44;
assign inst26_p17 = inst1_p46;
assign inst26_p20 = inst1_p49;
assign inst26_p21 = inst1_p50;
assign inst26_p23 = inst1_p52;
assign inst26_clk = clk;
assign inst26_p11 = inst1_p40;
assign inst26_p25 = inst1_p54;
assign inst26_p36 = inst1_p65;
assign inst26_p5 = inst1_p34;
assign inst26_p8 = inst1_p37;
assign inst26_p10 = inst1_p39;
assign inst26_reset = reset;
assign inst26_p13 = inst1_p42;
assign inst26_p18 = inst1_p47;
assign inst26_p30 = inst1_p59;
assign inst26_p7 = inst1_p36;
assign inst26_p24 = inst1_p53;
assign inst26_p32 = inst1_p61;
assign inst26_p14 = inst1_p43;
assign inst26_p26 = inst1_p55;
assign inst26_p31 = inst1_p60;
assign inst26_p27 = inst1_p56;
assign inst26_p33 = inst1_p62;
assign inst26_p22 = inst1_p51;
assign inst26_p34 = inst1_p63;
assign inst26_p35 = inst1_p64;
assign inst2_clk = clk;
assign inst2_reset = reset;
assign inst4_clk = clk;
assign inst4_reset = reset;
assign inst4_in =
  _guard2863 ? inst32_p37 :
  _guard2866 ? inst28_p37 :
  _guard2869 ? inst30_p37 :
  _guard2872 ? inst26_p37 :
  'x;
assign inst10_p4 = inst9_out;
assign inst10_clk = clk;
assign inst10_reset = reset;
assign inst11_p19 = inst3_p48;
assign inst11_p28 = inst3_p57;
assign inst11_p29 = inst3_p58;
assign inst11_p12 = inst3_p41;
assign inst11_p16 = inst3_p45;
assign inst11_p6 = inst3_p35;
assign inst11_p9 = inst3_p38;
assign inst11_p15 = inst3_p44;
assign inst11_p17 = inst3_p46;
assign inst11_p20 = inst3_p49;
assign inst11_p21 = inst3_p50;
assign inst11_p23 = inst3_p52;
assign inst11_clk = clk;
assign inst11_p11 = inst3_p40;
assign inst11_p25 = inst3_p54;
assign inst11_p36 = inst3_p65;
assign inst11_p5 = inst3_p34;
assign inst11_p8 = inst3_p37;
assign inst11_p10 = inst3_p39;
assign inst11_reset = reset;
assign inst11_p13 = inst3_p42;
assign inst11_p18 = inst3_p47;
assign inst11_p30 = inst3_p59;
assign inst11_p7 = inst3_p36;
assign inst11_p24 = inst3_p53;
assign inst11_p32 = inst3_p61;
assign inst11_p14 = inst3_p43;
assign inst11_p26 = inst3_p55;
assign inst11_p31 = inst3_p60;
assign inst11_p27 = inst3_p56;
assign inst11_p33 = inst3_p62;
assign inst11_p22 = inst3_p51;
assign inst11_p34 = inst3_p63;
assign inst11_p35 = inst3_p64;
assign inst13_p4 = inst9_out;
assign inst13_clk = clk;
assign inst13_reset = reset;
// COMPONENT END: comp92
endmodule
module comp93(
  input logic [31:0] p8,
  input logic [31:0] p9,
  input logic [31:0] p10,
  input logic [31:0] p11,
  input logic [31:0] p12,
  input logic [31:0] p13,
  input logic [31:0] p14,
  input logic [31:0] p15,
  input logic [31:0] p16,
  input logic [31:0] p17,
  input logic [31:0] p18,
  input logic [31:0] p19,
  input logic [31:0] p20,
  input logic [31:0] p21,
  input logic [31:0] p22,
  input logic [31:0] p23,
  input logic [31:0] p24,
  input logic [31:0] p25,
  input logic [31:0] p26,
  input logic [31:0] p27,
  input logic [31:0] p28,
  input logic [31:0] p29,
  input logic [31:0] p30,
  input logic [31:0] p31,
  input logic [31:0] p32,
  input logic [31:0] p33,
  input logic [31:0] p34,
  input logic [31:0] p35,
  input logic [31:0] p36,
  input logic [31:0] p37,
  input logic [31:0] p38,
  input logic [31:0] p39,
  output logic [1023:0] p40,
  input logic ev0,
  input logic clk,
  input logic reset
);
// COMPONENT START: comp93
logic [6:0] ev00__0state;
logic ev00__0_0;
logic [6:0] ev00__1state;
logic ev00__1_0;
logic ev00_clk;
logic ev00_reset;
logic ev00_go;
logic ev00_done;
logic [31:0] inst0_p108;
logic [31:0] inst0_p109;
logic [31:0] inst0_p110;
logic [31:0] inst0_p111;
logic [31:0] inst0_p112;
logic [31:0] inst0_p113;
logic [31:0] inst0_p114;
logic [31:0] inst0_p115;
logic [31:0] inst0_p116;
logic [31:0] inst0_p117;
logic [31:0] inst0_p118;
logic [31:0] inst0_p119;
logic [31:0] inst0_p120;
logic [31:0] inst0_p121;
logic [31:0] inst0_p122;
logic [31:0] inst0_p123;
logic [31:0] inst0_p124;
logic [31:0] inst0_p125;
logic [31:0] inst0_p126;
logic [31:0] inst0_p127;
logic [31:0] inst0_p128;
logic [31:0] inst0_p129;
logic [31:0] inst0_p130;
logic [31:0] inst0_p131;
logic [31:0] inst0_p132;
logic [31:0] inst0_p133;
logic [31:0] inst0_p134;
logic [31:0] inst0_p135;
logic [31:0] inst0_p136;
logic [31:0] inst0_p137;
logic [31:0] inst0_p138;
logic [31:0] inst0_p139;
logic [31:0] inst0_p140;
logic [31:0] inst0_p141;
logic [31:0] inst0_p142;
logic [31:0] inst0_p143;
logic [31:0] inst0_p144;
logic [31:0] inst0_p145;
logic [31:0] inst0_p146;
logic [31:0] inst0_p147;
logic [31:0] inst0_p148;
logic [31:0] inst0_p149;
logic [31:0] inst0_p150;
logic [31:0] inst0_p151;
logic [31:0] inst0_p152;
logic [31:0] inst0_p153;
logic [31:0] inst0_p154;
logic [31:0] inst0_p155;
logic [31:0] inst0_p156;
logic [31:0] inst0_p157;
logic [31:0] inst0_p158;
logic [31:0] inst0_p159;
logic [31:0] inst0_p160;
logic [31:0] inst0_p161;
logic [31:0] inst0_p162;
logic [31:0] inst0_p163;
logic [31:0] inst0_p164;
logic [31:0] inst0_p165;
logic [31:0] inst0_p166;
logic [31:0] inst0_p167;
logic [31:0] inst0_p168;
logic [31:0] inst0_p169;
logic [31:0] inst0_p170;
logic [31:0] inst0_p171;
logic inst0_ev0;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_p7;
logic [31:0] inst1_p8;
logic [31:0] inst1_p9;
logic [31:0] inst1_p10;
logic [31:0] inst1_p11;
logic [31:0] inst1_p12;
logic [31:0] inst1_p13;
logic [31:0] inst1_p14;
logic [31:0] inst1_p15;
logic [31:0] inst1_p16;
logic [31:0] inst1_p17;
logic [31:0] inst1_p18;
logic [31:0] inst1_p19;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic [31:0] inst1_p30;
logic [31:0] inst1_p31;
logic [31:0] inst1_p32;
logic [31:0] inst1_p33;
logic [31:0] inst1_p34;
logic [31:0] inst1_p35;
logic [31:0] inst1_p36;
logic [31:0] inst1_p37;
logic [31:0] inst1_p38;
logic [1023:0] inst1_p39;
logic inst1_reset;
logic inst1_clk;
counter_chain_2_128 ev00 (
    ._0_0(ev00__0_0),
    ._0state(ev00__0state),
    ._1_0(ev00__1_0),
    ._1state(ev00__1state),
    .clk(ev00_clk),
    .done(ev00_done),
    .go(ev00_go),
    .reset(ev00_reset)
);
comp92 inst0 (
    .clk(inst0_clk),
    .ev0(inst0_ev0),
    .p108(inst0_p108),
    .p109(inst0_p109),
    .p110(inst0_p110),
    .p111(inst0_p111),
    .p112(inst0_p112),
    .p113(inst0_p113),
    .p114(inst0_p114),
    .p115(inst0_p115),
    .p116(inst0_p116),
    .p117(inst0_p117),
    .p118(inst0_p118),
    .p119(inst0_p119),
    .p120(inst0_p120),
    .p121(inst0_p121),
    .p122(inst0_p122),
    .p123(inst0_p123),
    .p124(inst0_p124),
    .p125(inst0_p125),
    .p126(inst0_p126),
    .p127(inst0_p127),
    .p128(inst0_p128),
    .p129(inst0_p129),
    .p130(inst0_p130),
    .p131(inst0_p131),
    .p132(inst0_p132),
    .p133(inst0_p133),
    .p134(inst0_p134),
    .p135(inst0_p135),
    .p136(inst0_p136),
    .p137(inst0_p137),
    .p138(inst0_p138),
    .p139(inst0_p139),
    .p140(inst0_p140),
    .p141(inst0_p141),
    .p142(inst0_p142),
    .p143(inst0_p143),
    .p144(inst0_p144),
    .p145(inst0_p145),
    .p146(inst0_p146),
    .p147(inst0_p147),
    .p148(inst0_p148),
    .p149(inst0_p149),
    .p150(inst0_p150),
    .p151(inst0_p151),
    .p152(inst0_p152),
    .p153(inst0_p153),
    .p154(inst0_p154),
    .p155(inst0_p155),
    .p156(inst0_p156),
    .p157(inst0_p157),
    .p158(inst0_p158),
    .p159(inst0_p159),
    .p160(inst0_p160),
    .p161(inst0_p161),
    .p162(inst0_p162),
    .p163(inst0_p163),
    .p164(inst0_p164),
    .p165(inst0_p165),
    .p166(inst0_p166),
    .p167(inst0_p167),
    .p168(inst0_p168),
    .p169(inst0_p169),
    .p170(inst0_p170),
    .p171(inst0_p171),
    .reset(inst0_reset)
);
comp90 inst1 (
    .clk(inst1_clk),
    .p10(inst1_p10),
    .p11(inst1_p11),
    .p12(inst1_p12),
    .p13(inst1_p13),
    .p14(inst1_p14),
    .p15(inst1_p15),
    .p16(inst1_p16),
    .p17(inst1_p17),
    .p18(inst1_p18),
    .p19(inst1_p19),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .p30(inst1_p30),
    .p31(inst1_p31),
    .p32(inst1_p32),
    .p33(inst1_p33),
    .p34(inst1_p34),
    .p35(inst1_p35),
    .p36(inst1_p36),
    .p37(inst1_p37),
    .p38(inst1_p38),
    .p39(inst1_p39),
    .p7(inst1_p7),
    .p8(inst1_p8),
    .p9(inst1_p9),
    .reset(inst1_reset)
);
wire _guard0 = 1;
wire _guard1 = ev00__1_0;
wire _guard2 = ev00__1state >= 7'd1;
wire _guard3 = ev00__1state <= 7'd0;
wire _guard4 = _guard2 & _guard3;
wire _guard5 = _guard1 | _guard4;
wire _guard6 = ev00__1_0;
wire _guard7 = ev00__1state >= 7'd1;
wire _guard8 = ev00__1state <= 7'd0;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = _guard6 | _guard9;
wire _guard11 = ev00__1_0;
wire _guard12 = ev00__1state >= 7'd1;
wire _guard13 = ev00__1state <= 7'd0;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = _guard11 | _guard14;
wire _guard16 = ev00__1_0;
wire _guard17 = ev00__1state >= 7'd1;
wire _guard18 = ev00__1state <= 7'd0;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = _guard16 | _guard19;
wire _guard21 = ev00__1_0;
wire _guard22 = ev00__1state >= 7'd1;
wire _guard23 = ev00__1state <= 7'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard21 | _guard24;
wire _guard26 = ev00__1_0;
wire _guard27 = ev00__1state >= 7'd1;
wire _guard28 = ev00__1state <= 7'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard26 | _guard29;
wire _guard31 = ev00__1_0;
wire _guard32 = ev00__1state >= 7'd1;
wire _guard33 = ev00__1state <= 7'd0;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = _guard31 | _guard34;
wire _guard36 = ev00__1_0;
wire _guard37 = ev00__1state >= 7'd1;
wire _guard38 = ev00__1state <= 7'd0;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = _guard36 | _guard39;
wire _guard41 = ev00__1_0;
wire _guard42 = ev00__1state >= 7'd1;
wire _guard43 = ev00__1state <= 7'd0;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = _guard41 | _guard44;
wire _guard46 = ev00__1_0;
wire _guard47 = ev00__1state >= 7'd1;
wire _guard48 = ev00__1state <= 7'd0;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = _guard46 | _guard49;
wire _guard51 = ev00__1_0;
wire _guard52 = ev00__1state >= 7'd1;
wire _guard53 = ev00__1state <= 7'd0;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = _guard51 | _guard54;
wire _guard56 = ev00__1_0;
wire _guard57 = ev00__1state >= 7'd1;
wire _guard58 = ev00__1state <= 7'd0;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = _guard56 | _guard59;
wire _guard61 = ev00__1_0;
wire _guard62 = ev00__1state >= 7'd1;
wire _guard63 = ev00__1state <= 7'd0;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = _guard61 | _guard64;
wire _guard66 = ev00__1_0;
wire _guard67 = ev00__1state >= 7'd1;
wire _guard68 = ev00__1state <= 7'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = _guard66 | _guard69;
wire _guard71 = ev00__1_0;
wire _guard72 = ev00__1state >= 7'd1;
wire _guard73 = ev00__1state <= 7'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard71 | _guard74;
wire _guard76 = ev00__1_0;
wire _guard77 = ev00__1state >= 7'd1;
wire _guard78 = ev00__1state <= 7'd0;
wire _guard79 = _guard77 & _guard78;
wire _guard80 = _guard76 | _guard79;
wire _guard81 = ev00__1_0;
wire _guard82 = ev00__1state >= 7'd1;
wire _guard83 = ev00__1state <= 7'd0;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = _guard81 | _guard84;
wire _guard86 = ev00__1_0;
wire _guard87 = ev00__1state >= 7'd1;
wire _guard88 = ev00__1state <= 7'd0;
wire _guard89 = _guard87 & _guard88;
wire _guard90 = _guard86 | _guard89;
wire _guard91 = ev00__1_0;
wire _guard92 = ev00__1state >= 7'd1;
wire _guard93 = ev00__1state <= 7'd0;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = _guard91 | _guard94;
wire _guard96 = ev00__1_0;
wire _guard97 = ev00__1state >= 7'd1;
wire _guard98 = ev00__1state <= 7'd0;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = _guard96 | _guard99;
wire _guard101 = ev00__1_0;
wire _guard102 = ev00__1state >= 7'd1;
wire _guard103 = ev00__1state <= 7'd0;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = _guard101 | _guard104;
wire _guard106 = ev00__1_0;
wire _guard107 = ev00__1state >= 7'd1;
wire _guard108 = ev00__1state <= 7'd0;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = _guard106 | _guard109;
wire _guard111 = ev00__1_0;
wire _guard112 = ev00__1state >= 7'd1;
wire _guard113 = ev00__1state <= 7'd0;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = _guard111 | _guard114;
wire _guard116 = ev00__1_0;
wire _guard117 = ev00__1state >= 7'd1;
wire _guard118 = ev00__1state <= 7'd0;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = _guard116 | _guard119;
wire _guard121 = ev00__1_0;
wire _guard122 = ev00__1state >= 7'd1;
wire _guard123 = ev00__1state <= 7'd0;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = _guard121 | _guard124;
wire _guard126 = ev00__1_0;
wire _guard127 = ev00__1state >= 7'd1;
wire _guard128 = ev00__1state <= 7'd0;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = _guard126 | _guard129;
wire _guard131 = ev00__1_0;
wire _guard132 = ev00__1state >= 7'd1;
wire _guard133 = ev00__1state <= 7'd0;
wire _guard134 = _guard132 & _guard133;
wire _guard135 = _guard131 | _guard134;
wire _guard136 = ev00__1_0;
wire _guard137 = ev00__1state >= 7'd1;
wire _guard138 = ev00__1state <= 7'd0;
wire _guard139 = _guard137 & _guard138;
wire _guard140 = _guard136 | _guard139;
wire _guard141 = ev00__1_0;
wire _guard142 = ev00__1state >= 7'd1;
wire _guard143 = ev00__1state <= 7'd0;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = _guard141 | _guard144;
wire _guard146 = ev00__1_0;
wire _guard147 = ev00__1state >= 7'd1;
wire _guard148 = ev00__1state <= 7'd0;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = _guard146 | _guard149;
wire _guard151 = ev00__1_0;
wire _guard152 = ev00__1state >= 7'd1;
wire _guard153 = ev00__1state <= 7'd0;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = _guard151 | _guard154;
wire _guard156 = ev00__1_0;
wire _guard157 = ev00__1state >= 7'd1;
wire _guard158 = ev00__1state <= 7'd0;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = _guard156 | _guard159;
wire _guard161 = ev00__1_0;
wire _guard162 = ev00__1state >= 7'd1;
wire _guard163 = ev00__1state <= 7'd0;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = _guard161 | _guard164;
wire _guard166 = ev00__0_0;
wire _guard167 = ev00__0state >= 7'd1;
wire _guard168 = ev00__0state <= 7'd0;
wire _guard169 = _guard167 & _guard168;
wire _guard170 = _guard166 | _guard169;
wire _guard171 = ev00__0_0;
wire _guard172 = ev00__0state >= 7'd1;
wire _guard173 = ev00__0state <= 7'd0;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = _guard171 | _guard174;
wire _guard176 = ev00__0_0;
wire _guard177 = ev00__0state >= 7'd1;
wire _guard178 = ev00__0state <= 7'd0;
wire _guard179 = _guard177 & _guard178;
wire _guard180 = _guard176 | _guard179;
wire _guard181 = ev00__0_0;
wire _guard182 = ev00__0state >= 7'd1;
wire _guard183 = ev00__0state <= 7'd0;
wire _guard184 = _guard182 & _guard183;
wire _guard185 = _guard181 | _guard184;
wire _guard186 = ev00__0_0;
wire _guard187 = ev00__0state >= 7'd1;
wire _guard188 = ev00__0state <= 7'd0;
wire _guard189 = _guard187 & _guard188;
wire _guard190 = _guard186 | _guard189;
wire _guard191 = ev00__0_0;
wire _guard192 = ev00__0state >= 7'd1;
wire _guard193 = ev00__0state <= 7'd0;
wire _guard194 = _guard192 & _guard193;
wire _guard195 = _guard191 | _guard194;
wire _guard196 = ev00__0_0;
wire _guard197 = ev00__0state >= 7'd1;
wire _guard198 = ev00__0state <= 7'd0;
wire _guard199 = _guard197 & _guard198;
wire _guard200 = _guard196 | _guard199;
wire _guard201 = ev00__0_0;
wire _guard202 = ev00__0state >= 7'd1;
wire _guard203 = ev00__0state <= 7'd0;
wire _guard204 = _guard202 & _guard203;
wire _guard205 = _guard201 | _guard204;
wire _guard206 = ev00__0_0;
wire _guard207 = ev00__0state >= 7'd1;
wire _guard208 = ev00__0state <= 7'd0;
wire _guard209 = _guard207 & _guard208;
wire _guard210 = _guard206 | _guard209;
wire _guard211 = ev00__0_0;
wire _guard212 = ev00__0state >= 7'd1;
wire _guard213 = ev00__0state <= 7'd0;
wire _guard214 = _guard212 & _guard213;
wire _guard215 = _guard211 | _guard214;
wire _guard216 = ev00__0_0;
wire _guard217 = ev00__0state >= 7'd1;
wire _guard218 = ev00__0state <= 7'd0;
wire _guard219 = _guard217 & _guard218;
wire _guard220 = _guard216 | _guard219;
wire _guard221 = ev00__0_0;
wire _guard222 = ev00__0state >= 7'd1;
wire _guard223 = ev00__0state <= 7'd0;
wire _guard224 = _guard222 & _guard223;
wire _guard225 = _guard221 | _guard224;
wire _guard226 = ev00__0_0;
wire _guard227 = ev00__0state >= 7'd1;
wire _guard228 = ev00__0state <= 7'd0;
wire _guard229 = _guard227 & _guard228;
wire _guard230 = _guard226 | _guard229;
wire _guard231 = ev00__0_0;
wire _guard232 = ev00__0state >= 7'd1;
wire _guard233 = ev00__0state <= 7'd0;
wire _guard234 = _guard232 & _guard233;
wire _guard235 = _guard231 | _guard234;
wire _guard236 = ev00__0_0;
wire _guard237 = ev00__0state >= 7'd1;
wire _guard238 = ev00__0state <= 7'd0;
wire _guard239 = _guard237 & _guard238;
wire _guard240 = _guard236 | _guard239;
wire _guard241 = ev00__0_0;
wire _guard242 = ev00__0state >= 7'd1;
wire _guard243 = ev00__0state <= 7'd0;
wire _guard244 = _guard242 & _guard243;
wire _guard245 = _guard241 | _guard244;
wire _guard246 = ev00__0_0;
wire _guard247 = ev00__0state >= 7'd1;
wire _guard248 = ev00__0state <= 7'd0;
wire _guard249 = _guard247 & _guard248;
wire _guard250 = _guard246 | _guard249;
wire _guard251 = ev00__0_0;
wire _guard252 = ev00__0state >= 7'd1;
wire _guard253 = ev00__0state <= 7'd0;
wire _guard254 = _guard252 & _guard253;
wire _guard255 = _guard251 | _guard254;
wire _guard256 = ev00__0_0;
wire _guard257 = ev00__0state >= 7'd1;
wire _guard258 = ev00__0state <= 7'd0;
wire _guard259 = _guard257 & _guard258;
wire _guard260 = _guard256 | _guard259;
wire _guard261 = ev00__0_0;
wire _guard262 = ev00__0state >= 7'd1;
wire _guard263 = ev00__0state <= 7'd0;
wire _guard264 = _guard262 & _guard263;
wire _guard265 = _guard261 | _guard264;
wire _guard266 = ev00__0_0;
wire _guard267 = ev00__0state >= 7'd1;
wire _guard268 = ev00__0state <= 7'd0;
wire _guard269 = _guard267 & _guard268;
wire _guard270 = _guard266 | _guard269;
wire _guard271 = ev00__0_0;
wire _guard272 = ev00__0state >= 7'd1;
wire _guard273 = ev00__0state <= 7'd0;
wire _guard274 = _guard272 & _guard273;
wire _guard275 = _guard271 | _guard274;
wire _guard276 = ev00__0_0;
wire _guard277 = ev00__0state >= 7'd1;
wire _guard278 = ev00__0state <= 7'd0;
wire _guard279 = _guard277 & _guard278;
wire _guard280 = _guard276 | _guard279;
wire _guard281 = ev00__0_0;
wire _guard282 = ev00__0state >= 7'd1;
wire _guard283 = ev00__0state <= 7'd0;
wire _guard284 = _guard282 & _guard283;
wire _guard285 = _guard281 | _guard284;
wire _guard286 = ev00__0_0;
wire _guard287 = ev00__0state >= 7'd1;
wire _guard288 = ev00__0state <= 7'd0;
wire _guard289 = _guard287 & _guard288;
wire _guard290 = _guard286 | _guard289;
wire _guard291 = ev00__0_0;
wire _guard292 = ev00__0state >= 7'd1;
wire _guard293 = ev00__0state <= 7'd0;
wire _guard294 = _guard292 & _guard293;
wire _guard295 = _guard291 | _guard294;
wire _guard296 = ev00__0_0;
wire _guard297 = ev00__0state >= 7'd1;
wire _guard298 = ev00__0state <= 7'd0;
wire _guard299 = _guard297 & _guard298;
wire _guard300 = _guard296 | _guard299;
wire _guard301 = ev00__0_0;
wire _guard302 = ev00__0state >= 7'd1;
wire _guard303 = ev00__0state <= 7'd0;
wire _guard304 = _guard302 & _guard303;
wire _guard305 = _guard301 | _guard304;
wire _guard306 = ev00__0_0;
wire _guard307 = ev00__0state >= 7'd1;
wire _guard308 = ev00__0state <= 7'd0;
wire _guard309 = _guard307 & _guard308;
wire _guard310 = _guard306 | _guard309;
wire _guard311 = ev00__0_0;
wire _guard312 = ev00__0state >= 7'd1;
wire _guard313 = ev00__0state <= 7'd0;
wire _guard314 = _guard312 & _guard313;
wire _guard315 = _guard311 | _guard314;
wire _guard316 = ev00__0_0;
wire _guard317 = ev00__0state >= 7'd1;
wire _guard318 = ev00__0state <= 7'd0;
wire _guard319 = _guard317 & _guard318;
wire _guard320 = _guard316 | _guard319;
wire _guard321 = ev00__0_0;
wire _guard322 = ev00__0state >= 7'd1;
wire _guard323 = ev00__0state <= 7'd0;
wire _guard324 = _guard322 & _guard323;
wire _guard325 = _guard321 | _guard324;
wire _guard326 = ev00__0_0;
wire _guard327 = ev00__0state >= 7'd1;
wire _guard328 = ev00__0state <= 7'd0;
wire _guard329 = _guard327 & _guard328;
wire _guard330 = _guard326 | _guard329;
assign p40 =
  _guard5 ? inst1_p39 :
  1024'd0;
assign inst1_p19 = inst0_p152;
assign inst1_p28 = inst0_p161;
assign inst1_p29 = inst0_p162;
assign inst1_p38 = inst0_p171;
assign inst1_p12 = inst0_p145;
assign inst1_p16 = inst0_p149;
assign inst1_p9 = inst0_p142;
assign inst1_p15 = inst0_p148;
assign inst1_p17 = inst0_p150;
assign inst1_p20 = inst0_p153;
assign inst1_p21 = inst0_p154;
assign inst1_p23 = inst0_p156;
assign inst1_clk = clk;
assign inst1_p11 = inst0_p144;
assign inst1_p25 = inst0_p158;
assign inst1_p36 = inst0_p169;
assign inst1_p8 = inst0_p141;
assign inst1_p10 = inst0_p143;
assign inst1_reset = reset;
assign inst1_p13 = inst0_p146;
assign inst1_p18 = inst0_p151;
assign inst1_p30 = inst0_p163;
assign inst1_p7 = inst0_p140;
assign inst1_p24 = inst0_p157;
assign inst1_p32 = inst0_p165;
assign inst1_p14 = inst0_p147;
assign inst1_p26 = inst0_p159;
assign inst1_p31 = inst0_p164;
assign inst1_p27 = inst0_p160;
assign inst1_p33 = inst0_p166;
assign inst1_p22 = inst0_p155;
assign inst1_p34 = inst0_p167;
assign inst1_p35 = inst0_p168;
assign inst1_p37 = inst0_p170;
assign inst0_p120 = p20;
assign inst0_p130 = p30;
assign inst0_p137 = p37;
assign inst0_p110 = p10;
assign inst0_p115 = p15;
assign inst0_p116 = p16;
assign inst0_ev0 = _guard200;
assign inst0_p126 = p26;
assign inst0_p129 = p29;
assign inst0_p121 = p21;
assign inst0_p131 = p31;
assign inst0_p109 = p9;
assign inst0_p111 = p11;
assign inst0_p139 = p39;
assign inst0_clk = clk;
assign inst0_p123 = p23;
assign inst0_p127 = p27;
assign inst0_p128 = p28;
assign inst0_p132 = p32;
assign inst0_p135 = p35;
assign inst0_p136 = p36;
assign inst0_reset = reset;
assign inst0_p113 = p13;
assign inst0_p117 = p17;
assign inst0_p133 = p33;
assign inst0_p119 = p19;
assign inst0_p112 = p12;
assign inst0_p108 = p8;
assign inst0_p125 = p25;
assign inst0_p114 = p14;
assign inst0_p118 = p18;
assign inst0_p138 = p38;
assign inst0_p122 = p22;
assign inst0_p124 = p24;
assign inst0_p134 = p34;
assign ev00_clk = clk;
assign ev00_go = ev0;
assign ev00_reset = reset;
// COMPONENT END: comp93
endmodule
module main(
  input logic [1023:0] in,
  output logic [1023:0] out,
  input logic go,
  input logic reset,
  input logic clk
);
// COMPONENT START: main
logic [6:0] go0__0state;
logic go0__0_0;
logic [6:0] go0__1state;
logic go0__1_0;
logic go0_clk;
logic go0_reset;
logic go0_go;
logic go0_done;
logic [1023:0] inst0_p8;
logic [31:0] inst0_p9;
logic [31:0] inst0_p10;
logic [31:0] inst0_p11;
logic [31:0] inst0_p12;
logic [31:0] inst0_p13;
logic [31:0] inst0_p14;
logic [31:0] inst0_p15;
logic [31:0] inst0_p16;
logic [31:0] inst0_p17;
logic [31:0] inst0_p18;
logic [31:0] inst0_p19;
logic [31:0] inst0_p20;
logic [31:0] inst0_p21;
logic [31:0] inst0_p22;
logic [31:0] inst0_p23;
logic [31:0] inst0_p24;
logic [31:0] inst0_p25;
logic [31:0] inst0_p26;
logic [31:0] inst0_p27;
logic [31:0] inst0_p28;
logic [31:0] inst0_p29;
logic [31:0] inst0_p30;
logic [31:0] inst0_p31;
logic [31:0] inst0_p32;
logic [31:0] inst0_p33;
logic [31:0] inst0_p34;
logic [31:0] inst0_p35;
logic [31:0] inst0_p36;
logic [31:0] inst0_p37;
logic [31:0] inst0_p38;
logic [31:0] inst0_p39;
logic [31:0] inst0_p40;
logic inst0_clk;
logic inst0_reset;
logic [31:0] inst1_p8;
logic [31:0] inst1_p9;
logic [31:0] inst1_p10;
logic [31:0] inst1_p11;
logic [31:0] inst1_p12;
logic [31:0] inst1_p13;
logic [31:0] inst1_p14;
logic [31:0] inst1_p15;
logic [31:0] inst1_p16;
logic [31:0] inst1_p17;
logic [31:0] inst1_p18;
logic [31:0] inst1_p19;
logic [31:0] inst1_p20;
logic [31:0] inst1_p21;
logic [31:0] inst1_p22;
logic [31:0] inst1_p23;
logic [31:0] inst1_p24;
logic [31:0] inst1_p25;
logic [31:0] inst1_p26;
logic [31:0] inst1_p27;
logic [31:0] inst1_p28;
logic [31:0] inst1_p29;
logic [31:0] inst1_p30;
logic [31:0] inst1_p31;
logic [31:0] inst1_p32;
logic [31:0] inst1_p33;
logic [31:0] inst1_p34;
logic [31:0] inst1_p35;
logic [31:0] inst1_p36;
logic [31:0] inst1_p37;
logic [31:0] inst1_p38;
logic [31:0] inst1_p39;
logic [1023:0] inst1_p40;
logic inst1_ev0;
logic inst1_clk;
logic inst1_reset;
counter_chain_2_128 go0 (
    ._0_0(go0__0_0),
    ._0state(go0__0state),
    ._1_0(go0__1_0),
    ._1state(go0__1state),
    .clk(go0_clk),
    .done(go0_done),
    .go(go0_go),
    .reset(go0_reset)
);
comp32 inst0 (
    .clk(inst0_clk),
    .p10(inst0_p10),
    .p11(inst0_p11),
    .p12(inst0_p12),
    .p13(inst0_p13),
    .p14(inst0_p14),
    .p15(inst0_p15),
    .p16(inst0_p16),
    .p17(inst0_p17),
    .p18(inst0_p18),
    .p19(inst0_p19),
    .p20(inst0_p20),
    .p21(inst0_p21),
    .p22(inst0_p22),
    .p23(inst0_p23),
    .p24(inst0_p24),
    .p25(inst0_p25),
    .p26(inst0_p26),
    .p27(inst0_p27),
    .p28(inst0_p28),
    .p29(inst0_p29),
    .p30(inst0_p30),
    .p31(inst0_p31),
    .p32(inst0_p32),
    .p33(inst0_p33),
    .p34(inst0_p34),
    .p35(inst0_p35),
    .p36(inst0_p36),
    .p37(inst0_p37),
    .p38(inst0_p38),
    .p39(inst0_p39),
    .p40(inst0_p40),
    .p8(inst0_p8),
    .p9(inst0_p9),
    .reset(inst0_reset)
);
comp93 inst1 (
    .clk(inst1_clk),
    .ev0(inst1_ev0),
    .p10(inst1_p10),
    .p11(inst1_p11),
    .p12(inst1_p12),
    .p13(inst1_p13),
    .p14(inst1_p14),
    .p15(inst1_p15),
    .p16(inst1_p16),
    .p17(inst1_p17),
    .p18(inst1_p18),
    .p19(inst1_p19),
    .p20(inst1_p20),
    .p21(inst1_p21),
    .p22(inst1_p22),
    .p23(inst1_p23),
    .p24(inst1_p24),
    .p25(inst1_p25),
    .p26(inst1_p26),
    .p27(inst1_p27),
    .p28(inst1_p28),
    .p29(inst1_p29),
    .p30(inst1_p30),
    .p31(inst1_p31),
    .p32(inst1_p32),
    .p33(inst1_p33),
    .p34(inst1_p34),
    .p35(inst1_p35),
    .p36(inst1_p36),
    .p37(inst1_p37),
    .p38(inst1_p38),
    .p39(inst1_p39),
    .p40(inst1_p40),
    .p8(inst1_p8),
    .p9(inst1_p9),
    .reset(inst1_reset)
);
wire _guard0 = 1;
wire _guard1 = go0__1_0;
wire _guard2 = go0__1state >= 7'd1;
wire _guard3 = go0__1state <= 7'd0;
wire _guard4 = _guard2 & _guard3;
wire _guard5 = _guard1 | _guard4;
wire _guard6 = go0__0_0;
wire _guard7 = go0__0state >= 7'd1;
wire _guard8 = go0__0state <= 7'd0;
wire _guard9 = _guard7 & _guard8;
wire _guard10 = _guard6 | _guard9;
wire _guard11 = go0__0_0;
wire _guard12 = go0__0state >= 7'd1;
wire _guard13 = go0__0state <= 7'd0;
wire _guard14 = _guard12 & _guard13;
wire _guard15 = _guard11 | _guard14;
wire _guard16 = go0__0_0;
wire _guard17 = go0__0state >= 7'd1;
wire _guard18 = go0__0state <= 7'd0;
wire _guard19 = _guard17 & _guard18;
wire _guard20 = _guard16 | _guard19;
wire _guard21 = go0__0_0;
wire _guard22 = go0__0state >= 7'd1;
wire _guard23 = go0__0state <= 7'd0;
wire _guard24 = _guard22 & _guard23;
wire _guard25 = _guard21 | _guard24;
wire _guard26 = go0__0_0;
wire _guard27 = go0__0state >= 7'd1;
wire _guard28 = go0__0state <= 7'd0;
wire _guard29 = _guard27 & _guard28;
wire _guard30 = _guard26 | _guard29;
wire _guard31 = go0__0_0;
wire _guard32 = go0__0state >= 7'd1;
wire _guard33 = go0__0state <= 7'd0;
wire _guard34 = _guard32 & _guard33;
wire _guard35 = _guard31 | _guard34;
wire _guard36 = go0__0_0;
wire _guard37 = go0__0state >= 7'd1;
wire _guard38 = go0__0state <= 7'd0;
wire _guard39 = _guard37 & _guard38;
wire _guard40 = _guard36 | _guard39;
wire _guard41 = go0__0_0;
wire _guard42 = go0__0state >= 7'd1;
wire _guard43 = go0__0state <= 7'd0;
wire _guard44 = _guard42 & _guard43;
wire _guard45 = _guard41 | _guard44;
wire _guard46 = go0__0_0;
wire _guard47 = go0__0state >= 7'd1;
wire _guard48 = go0__0state <= 7'd0;
wire _guard49 = _guard47 & _guard48;
wire _guard50 = _guard46 | _guard49;
wire _guard51 = go0__0_0;
wire _guard52 = go0__0state >= 7'd1;
wire _guard53 = go0__0state <= 7'd0;
wire _guard54 = _guard52 & _guard53;
wire _guard55 = _guard51 | _guard54;
wire _guard56 = go0__0_0;
wire _guard57 = go0__0state >= 7'd1;
wire _guard58 = go0__0state <= 7'd0;
wire _guard59 = _guard57 & _guard58;
wire _guard60 = _guard56 | _guard59;
wire _guard61 = go0__0_0;
wire _guard62 = go0__0state >= 7'd1;
wire _guard63 = go0__0state <= 7'd0;
wire _guard64 = _guard62 & _guard63;
wire _guard65 = _guard61 | _guard64;
wire _guard66 = go0__0_0;
wire _guard67 = go0__0state >= 7'd1;
wire _guard68 = go0__0state <= 7'd0;
wire _guard69 = _guard67 & _guard68;
wire _guard70 = _guard66 | _guard69;
wire _guard71 = go0__0_0;
wire _guard72 = go0__0state >= 7'd1;
wire _guard73 = go0__0state <= 7'd0;
wire _guard74 = _guard72 & _guard73;
wire _guard75 = _guard71 | _guard74;
wire _guard76 = go0__0_0;
wire _guard77 = go0__0state >= 7'd1;
wire _guard78 = go0__0state <= 7'd0;
wire _guard79 = _guard77 & _guard78;
wire _guard80 = _guard76 | _guard79;
wire _guard81 = go0__0_0;
wire _guard82 = go0__0state >= 7'd1;
wire _guard83 = go0__0state <= 7'd0;
wire _guard84 = _guard82 & _guard83;
wire _guard85 = _guard81 | _guard84;
wire _guard86 = go0__0_0;
wire _guard87 = go0__0state >= 7'd1;
wire _guard88 = go0__0state <= 7'd0;
wire _guard89 = _guard87 & _guard88;
wire _guard90 = _guard86 | _guard89;
wire _guard91 = go0__0_0;
wire _guard92 = go0__0state >= 7'd1;
wire _guard93 = go0__0state <= 7'd0;
wire _guard94 = _guard92 & _guard93;
wire _guard95 = _guard91 | _guard94;
wire _guard96 = go0__0_0;
wire _guard97 = go0__0state >= 7'd1;
wire _guard98 = go0__0state <= 7'd0;
wire _guard99 = _guard97 & _guard98;
wire _guard100 = _guard96 | _guard99;
wire _guard101 = go0__0_0;
wire _guard102 = go0__0state >= 7'd1;
wire _guard103 = go0__0state <= 7'd0;
wire _guard104 = _guard102 & _guard103;
wire _guard105 = _guard101 | _guard104;
wire _guard106 = go0__0_0;
wire _guard107 = go0__0state >= 7'd1;
wire _guard108 = go0__0state <= 7'd0;
wire _guard109 = _guard107 & _guard108;
wire _guard110 = _guard106 | _guard109;
wire _guard111 = go0__0_0;
wire _guard112 = go0__0state >= 7'd1;
wire _guard113 = go0__0state <= 7'd0;
wire _guard114 = _guard112 & _guard113;
wire _guard115 = _guard111 | _guard114;
wire _guard116 = go0__0_0;
wire _guard117 = go0__0state >= 7'd1;
wire _guard118 = go0__0state <= 7'd0;
wire _guard119 = _guard117 & _guard118;
wire _guard120 = _guard116 | _guard119;
wire _guard121 = go0__0_0;
wire _guard122 = go0__0state >= 7'd1;
wire _guard123 = go0__0state <= 7'd0;
wire _guard124 = _guard122 & _guard123;
wire _guard125 = _guard121 | _guard124;
wire _guard126 = go0__0_0;
wire _guard127 = go0__0state >= 7'd1;
wire _guard128 = go0__0state <= 7'd0;
wire _guard129 = _guard127 & _guard128;
wire _guard130 = _guard126 | _guard129;
wire _guard131 = go0__0_0;
wire _guard132 = go0__0state >= 7'd1;
wire _guard133 = go0__0state <= 7'd0;
wire _guard134 = _guard132 & _guard133;
wire _guard135 = _guard131 | _guard134;
wire _guard136 = go0__0_0;
wire _guard137 = go0__0state >= 7'd1;
wire _guard138 = go0__0state <= 7'd0;
wire _guard139 = _guard137 & _guard138;
wire _guard140 = _guard136 | _guard139;
wire _guard141 = go0__0_0;
wire _guard142 = go0__0state >= 7'd1;
wire _guard143 = go0__0state <= 7'd0;
wire _guard144 = _guard142 & _guard143;
wire _guard145 = _guard141 | _guard144;
wire _guard146 = go0__0_0;
wire _guard147 = go0__0state >= 7'd1;
wire _guard148 = go0__0state <= 7'd0;
wire _guard149 = _guard147 & _guard148;
wire _guard150 = _guard146 | _guard149;
wire _guard151 = go0__0_0;
wire _guard152 = go0__0state >= 7'd1;
wire _guard153 = go0__0state <= 7'd0;
wire _guard154 = _guard152 & _guard153;
wire _guard155 = _guard151 | _guard154;
wire _guard156 = go0__0_0;
wire _guard157 = go0__0state >= 7'd1;
wire _guard158 = go0__0state <= 7'd0;
wire _guard159 = _guard157 & _guard158;
wire _guard160 = _guard156 | _guard159;
wire _guard161 = go0__0_0;
wire _guard162 = go0__0state >= 7'd1;
wire _guard163 = go0__0state <= 7'd0;
wire _guard164 = _guard162 & _guard163;
wire _guard165 = _guard161 | _guard164;
wire _guard166 = go0__0_0;
wire _guard167 = go0__0state >= 7'd1;
wire _guard168 = go0__0state <= 7'd0;
wire _guard169 = _guard167 & _guard168;
wire _guard170 = _guard166 | _guard169;
wire _guard171 = go0__0_0;
wire _guard172 = go0__0state >= 7'd1;
wire _guard173 = go0__0state <= 7'd0;
wire _guard174 = _guard172 & _guard173;
wire _guard175 = _guard171 | _guard174;
assign out =
  _guard5 ? inst1_p40 :
  1024'd0;
assign go0_clk = clk;
assign go0_go = go;
assign go0_reset = reset;
assign inst1_p19 = inst0_p20;
assign inst1_p28 = inst0_p29;
assign inst1_p29 = inst0_p30;
assign inst1_p38 = inst0_p39;
assign inst1_p12 = inst0_p13;
assign inst1_p16 = inst0_p17;
assign inst1_ev0 = _guard40;
assign inst1_p9 = inst0_p10;
assign inst1_p15 = inst0_p16;
assign inst1_p17 = inst0_p18;
assign inst1_p20 = inst0_p21;
assign inst1_p21 = inst0_p22;
assign inst1_p23 = inst0_p24;
assign inst1_clk = clk;
assign inst1_p11 = inst0_p12;
assign inst1_p25 = inst0_p26;
assign inst1_p36 = inst0_p37;
assign inst1_p39 = inst0_p40;
assign inst1_p8 = inst0_p9;
assign inst1_p10 = inst0_p11;
assign inst1_reset = reset;
assign inst1_p13 = inst0_p14;
assign inst1_p18 = inst0_p19;
assign inst1_p30 = inst0_p31;
assign inst1_p24 = inst0_p25;
assign inst1_p32 = inst0_p33;
assign inst1_p14 = inst0_p15;
assign inst1_p26 = inst0_p27;
assign inst1_p31 = inst0_p32;
assign inst1_p27 = inst0_p28;
assign inst1_p33 = inst0_p34;
assign inst1_p22 = inst0_p23;
assign inst1_p34 = inst0_p35;
assign inst1_p35 = inst0_p36;
assign inst1_p37 = inst0_p38;
assign inst0_clk = clk;
assign inst0_p8 = in;
assign inst0_reset = reset;
// COMPONENT END: main
endmodule
module counter_chain_2_128(
  output logic [6:0] _0state,
  output logic _0_0,
  output logic [6:0] _1state,
  output logic _1_0,
  input logic clk,
  input logic reset,
  input logic go,
  output logic done
);
// COMPONENT START: counter_chain_2_128
logic c0_clk;
logic c0_reset;
logic [6:0] c0_state;
logic c0__0;
logic c0_go;
logic c0_done;
logic c1_clk;
logic c1_reset;
logic [6:0] c1_state;
logic c1__0;
logic c1_go;
logic c1_done;
counter_128 c0 (
    ._0(c0__0),
    .clk(c0_clk),
    .done(c0_done),
    .go(c0_go),
    .reset(c0_reset),
    .state(c0_state)
);
counter_128 c1 (
    ._0(c1__0),
    .clk(c1_clk),
    .done(c1_done),
    .go(c1_go),
    .reset(c1_reset),
    .state(c1_state)
);
wire _guard0 = 1;
assign done = c1_done;
assign _0state = c0_state;
assign _1state = c1_state;
assign _0_0 = c0__0;
assign _1_0 = c1__0;
assign c1_clk = clk;
assign c1_go = c0_done;
assign c1_reset = reset;
assign c0_clk = clk;
assign c0_go = go;
assign c0_reset = reset;
// COMPONENT END: counter_chain_2_128
endmodule
module fsm_31(
  output logic _0,
  output logic _1,
  output logic _2,
  output logic _3,
  output logic _4,
  output logic _5,
  output logic _6,
  output logic _7,
  output logic _8,
  output logic _9,
  output logic _10,
  output logic _11,
  output logic _12,
  output logic _13,
  output logic _14,
  output logic _15,
  output logic _16,
  output logic _17,
  output logic _18,
  output logic _19,
  output logic _20,
  output logic _21,
  output logic _22,
  output logic _23,
  output logic _24,
  output logic _25,
  output logic _26,
  output logic _27,
  output logic _28,
  output logic _29,
  output logic _30,
  input logic clk,
  input logic reset,
  input logic go,
  output logic done
);
// COMPONENT START: fsm_31
logic r_in;
logic r_write_en;
logic r_clk;
logic r_reset;
logic r_out;
logic r_done;
logic r0_in;
logic r0_write_en;
logic r0_clk;
logic r0_reset;
logic r0_out;
logic r0_done;
logic r1_in;
logic r1_write_en;
logic r1_clk;
logic r1_reset;
logic r1_out;
logic r1_done;
logic r2_in;
logic r2_write_en;
logic r2_clk;
logic r2_reset;
logic r2_out;
logic r2_done;
logic r3_in;
logic r3_write_en;
logic r3_clk;
logic r3_reset;
logic r3_out;
logic r3_done;
logic r4_in;
logic r4_write_en;
logic r4_clk;
logic r4_reset;
logic r4_out;
logic r4_done;
logic r5_in;
logic r5_write_en;
logic r5_clk;
logic r5_reset;
logic r5_out;
logic r5_done;
logic r6_in;
logic r6_write_en;
logic r6_clk;
logic r6_reset;
logic r6_out;
logic r6_done;
logic r7_in;
logic r7_write_en;
logic r7_clk;
logic r7_reset;
logic r7_out;
logic r7_done;
logic r8_in;
logic r8_write_en;
logic r8_clk;
logic r8_reset;
logic r8_out;
logic r8_done;
logic r9_in;
logic r9_write_en;
logic r9_clk;
logic r9_reset;
logic r9_out;
logic r9_done;
logic r10_in;
logic r10_write_en;
logic r10_clk;
logic r10_reset;
logic r10_out;
logic r10_done;
logic r11_in;
logic r11_write_en;
logic r11_clk;
logic r11_reset;
logic r11_out;
logic r11_done;
logic r12_in;
logic r12_write_en;
logic r12_clk;
logic r12_reset;
logic r12_out;
logic r12_done;
logic r13_in;
logic r13_write_en;
logic r13_clk;
logic r13_reset;
logic r13_out;
logic r13_done;
logic r14_in;
logic r14_write_en;
logic r14_clk;
logic r14_reset;
logic r14_out;
logic r14_done;
logic r15_in;
logic r15_write_en;
logic r15_clk;
logic r15_reset;
logic r15_out;
logic r15_done;
logic r16_in;
logic r16_write_en;
logic r16_clk;
logic r16_reset;
logic r16_out;
logic r16_done;
logic r17_in;
logic r17_write_en;
logic r17_clk;
logic r17_reset;
logic r17_out;
logic r17_done;
logic r18_in;
logic r18_write_en;
logic r18_clk;
logic r18_reset;
logic r18_out;
logic r18_done;
logic r19_in;
logic r19_write_en;
logic r19_clk;
logic r19_reset;
logic r19_out;
logic r19_done;
logic r20_in;
logic r20_write_en;
logic r20_clk;
logic r20_reset;
logic r20_out;
logic r20_done;
logic r21_in;
logic r21_write_en;
logic r21_clk;
logic r21_reset;
logic r21_out;
logic r21_done;
logic r22_in;
logic r22_write_en;
logic r22_clk;
logic r22_reset;
logic r22_out;
logic r22_done;
logic r23_in;
logic r23_write_en;
logic r23_clk;
logic r23_reset;
logic r23_out;
logic r23_done;
logic r24_in;
logic r24_write_en;
logic r24_clk;
logic r24_reset;
logic r24_out;
logic r24_done;
logic r25_in;
logic r25_write_en;
logic r25_clk;
logic r25_reset;
logic r25_out;
logic r25_done;
logic r26_in;
logic r26_write_en;
logic r26_clk;
logic r26_reset;
logic r26_out;
logic r26_done;
logic r27_in;
logic r27_write_en;
logic r27_clk;
logic r27_reset;
logic r27_out;
logic r27_done;
logic r28_in;
logic r28_write_en;
logic r28_clk;
logic r28_reset;
logic r28_out;
logic r28_done;
logic r29_in;
logic r29_write_en;
logic r29_clk;
logic r29_reset;
logic r29_out;
logic r29_done;
std_reg # (
    .WIDTH(1)
) r (
    .clk(r_clk),
    .done(r_done),
    .in(r_in),
    .out(r_out),
    .reset(r_reset),
    .write_en(r_write_en)
);
std_reg # (
    .WIDTH(1)
) r0 (
    .clk(r0_clk),
    .done(r0_done),
    .in(r0_in),
    .out(r0_out),
    .reset(r0_reset),
    .write_en(r0_write_en)
);
std_reg # (
    .WIDTH(1)
) r1 (
    .clk(r1_clk),
    .done(r1_done),
    .in(r1_in),
    .out(r1_out),
    .reset(r1_reset),
    .write_en(r1_write_en)
);
std_reg # (
    .WIDTH(1)
) r2 (
    .clk(r2_clk),
    .done(r2_done),
    .in(r2_in),
    .out(r2_out),
    .reset(r2_reset),
    .write_en(r2_write_en)
);
std_reg # (
    .WIDTH(1)
) r3 (
    .clk(r3_clk),
    .done(r3_done),
    .in(r3_in),
    .out(r3_out),
    .reset(r3_reset),
    .write_en(r3_write_en)
);
std_reg # (
    .WIDTH(1)
) r4 (
    .clk(r4_clk),
    .done(r4_done),
    .in(r4_in),
    .out(r4_out),
    .reset(r4_reset),
    .write_en(r4_write_en)
);
std_reg # (
    .WIDTH(1)
) r5 (
    .clk(r5_clk),
    .done(r5_done),
    .in(r5_in),
    .out(r5_out),
    .reset(r5_reset),
    .write_en(r5_write_en)
);
std_reg # (
    .WIDTH(1)
) r6 (
    .clk(r6_clk),
    .done(r6_done),
    .in(r6_in),
    .out(r6_out),
    .reset(r6_reset),
    .write_en(r6_write_en)
);
std_reg # (
    .WIDTH(1)
) r7 (
    .clk(r7_clk),
    .done(r7_done),
    .in(r7_in),
    .out(r7_out),
    .reset(r7_reset),
    .write_en(r7_write_en)
);
std_reg # (
    .WIDTH(1)
) r8 (
    .clk(r8_clk),
    .done(r8_done),
    .in(r8_in),
    .out(r8_out),
    .reset(r8_reset),
    .write_en(r8_write_en)
);
std_reg # (
    .WIDTH(1)
) r9 (
    .clk(r9_clk),
    .done(r9_done),
    .in(r9_in),
    .out(r9_out),
    .reset(r9_reset),
    .write_en(r9_write_en)
);
std_reg # (
    .WIDTH(1)
) r10 (
    .clk(r10_clk),
    .done(r10_done),
    .in(r10_in),
    .out(r10_out),
    .reset(r10_reset),
    .write_en(r10_write_en)
);
std_reg # (
    .WIDTH(1)
) r11 (
    .clk(r11_clk),
    .done(r11_done),
    .in(r11_in),
    .out(r11_out),
    .reset(r11_reset),
    .write_en(r11_write_en)
);
std_reg # (
    .WIDTH(1)
) r12 (
    .clk(r12_clk),
    .done(r12_done),
    .in(r12_in),
    .out(r12_out),
    .reset(r12_reset),
    .write_en(r12_write_en)
);
std_reg # (
    .WIDTH(1)
) r13 (
    .clk(r13_clk),
    .done(r13_done),
    .in(r13_in),
    .out(r13_out),
    .reset(r13_reset),
    .write_en(r13_write_en)
);
std_reg # (
    .WIDTH(1)
) r14 (
    .clk(r14_clk),
    .done(r14_done),
    .in(r14_in),
    .out(r14_out),
    .reset(r14_reset),
    .write_en(r14_write_en)
);
std_reg # (
    .WIDTH(1)
) r15 (
    .clk(r15_clk),
    .done(r15_done),
    .in(r15_in),
    .out(r15_out),
    .reset(r15_reset),
    .write_en(r15_write_en)
);
std_reg # (
    .WIDTH(1)
) r16 (
    .clk(r16_clk),
    .done(r16_done),
    .in(r16_in),
    .out(r16_out),
    .reset(r16_reset),
    .write_en(r16_write_en)
);
std_reg # (
    .WIDTH(1)
) r17 (
    .clk(r17_clk),
    .done(r17_done),
    .in(r17_in),
    .out(r17_out),
    .reset(r17_reset),
    .write_en(r17_write_en)
);
std_reg # (
    .WIDTH(1)
) r18 (
    .clk(r18_clk),
    .done(r18_done),
    .in(r18_in),
    .out(r18_out),
    .reset(r18_reset),
    .write_en(r18_write_en)
);
std_reg # (
    .WIDTH(1)
) r19 (
    .clk(r19_clk),
    .done(r19_done),
    .in(r19_in),
    .out(r19_out),
    .reset(r19_reset),
    .write_en(r19_write_en)
);
std_reg # (
    .WIDTH(1)
) r20 (
    .clk(r20_clk),
    .done(r20_done),
    .in(r20_in),
    .out(r20_out),
    .reset(r20_reset),
    .write_en(r20_write_en)
);
std_reg # (
    .WIDTH(1)
) r21 (
    .clk(r21_clk),
    .done(r21_done),
    .in(r21_in),
    .out(r21_out),
    .reset(r21_reset),
    .write_en(r21_write_en)
);
std_reg # (
    .WIDTH(1)
) r22 (
    .clk(r22_clk),
    .done(r22_done),
    .in(r22_in),
    .out(r22_out),
    .reset(r22_reset),
    .write_en(r22_write_en)
);
std_reg # (
    .WIDTH(1)
) r23 (
    .clk(r23_clk),
    .done(r23_done),
    .in(r23_in),
    .out(r23_out),
    .reset(r23_reset),
    .write_en(r23_write_en)
);
std_reg # (
    .WIDTH(1)
) r24 (
    .clk(r24_clk),
    .done(r24_done),
    .in(r24_in),
    .out(r24_out),
    .reset(r24_reset),
    .write_en(r24_write_en)
);
std_reg # (
    .WIDTH(1)
) r25 (
    .clk(r25_clk),
    .done(r25_done),
    .in(r25_in),
    .out(r25_out),
    .reset(r25_reset),
    .write_en(r25_write_en)
);
std_reg # (
    .WIDTH(1)
) r26 (
    .clk(r26_clk),
    .done(r26_done),
    .in(r26_in),
    .out(r26_out),
    .reset(r26_reset),
    .write_en(r26_write_en)
);
std_reg # (
    .WIDTH(1)
) r27 (
    .clk(r27_clk),
    .done(r27_done),
    .in(r27_in),
    .out(r27_out),
    .reset(r27_reset),
    .write_en(r27_write_en)
);
std_reg # (
    .WIDTH(1)
) r28 (
    .clk(r28_clk),
    .done(r28_done),
    .in(r28_in),
    .out(r28_out),
    .reset(r28_reset),
    .write_en(r28_write_en)
);
std_reg # (
    .WIDTH(1)
) r29 (
    .clk(r29_clk),
    .done(r29_done),
    .in(r29_in),
    .out(r29_out),
    .reset(r29_reset),
    .write_en(r29_write_en)
);
wire _guard0 = 1;
assign r5_write_en = 1'd1;
assign r5_clk = clk;
assign r5_reset = reset;
assign r5_in = r4_out;
assign done = r29_out;
assign _29 = r27_out;
assign _19 = r17_out;
assign _21 = r19_out;
assign _24 = r22_out;
assign _7 = r5_out;
assign _10 = r8_out;
assign _27 = r25_out;
assign _9 = r7_out;
assign _11 = r9_out;
assign _22 = r20_out;
assign _5 = r3_out;
assign _18 = r16_out;
assign _26 = r24_out;
assign _28 = r26_out;
assign _2 = r0_out;
assign _12 = r10_out;
assign _25 = r23_out;
assign _1 = r_out;
assign _15 = r13_out;
assign _23 = r21_out;
assign _14 = r12_out;
assign _0 = go;
assign _16 = r14_out;
assign _30 = r28_out;
assign _6 = r4_out;
assign _3 = r1_out;
assign _4 = r2_out;
assign _20 = r18_out;
assign _13 = r11_out;
assign _8 = r6_out;
assign _17 = r15_out;
assign r11_write_en = 1'd1;
assign r11_clk = clk;
assign r11_reset = reset;
assign r11_in = r10_out;
assign r13_write_en = 1'd1;
assign r13_clk = clk;
assign r13_reset = reset;
assign r13_in = r12_out;
assign r18_write_en = 1'd1;
assign r18_clk = clk;
assign r18_reset = reset;
assign r18_in = r17_out;
assign r20_write_en = 1'd1;
assign r20_clk = clk;
assign r20_reset = reset;
assign r20_in = r19_out;
assign r26_write_en = 1'd1;
assign r26_clk = clk;
assign r26_reset = reset;
assign r26_in = r25_out;
assign r27_write_en = 1'd1;
assign r27_clk = clk;
assign r27_reset = reset;
assign r27_in = r26_out;
assign r25_write_en = 1'd1;
assign r25_clk = clk;
assign r25_reset = reset;
assign r25_in = r24_out;
assign r19_write_en = 1'd1;
assign r19_clk = clk;
assign r19_reset = reset;
assign r19_in = r18_out;
assign r10_write_en = 1'd1;
assign r10_clk = clk;
assign r10_reset = reset;
assign r10_in = r9_out;
assign r15_write_en = 1'd1;
assign r15_clk = clk;
assign r15_reset = reset;
assign r15_in = r14_out;
assign r22_write_en = 1'd1;
assign r22_clk = clk;
assign r22_reset = reset;
assign r22_in = r21_out;
assign r28_write_en = 1'd1;
assign r28_clk = clk;
assign r28_reset = reset;
assign r28_in = r27_out;
assign r12_write_en = 1'd1;
assign r12_clk = clk;
assign r12_reset = reset;
assign r12_in = r11_out;
assign r_write_en = 1'd1;
assign r_clk = clk;
assign r_reset = reset;
assign r_in = go;
assign r0_write_en = 1'd1;
assign r0_clk = clk;
assign r0_reset = reset;
assign r0_in = r_out;
assign r1_write_en = 1'd1;
assign r1_clk = clk;
assign r1_reset = reset;
assign r1_in = r0_out;
assign r23_write_en = 1'd1;
assign r23_clk = clk;
assign r23_reset = reset;
assign r23_in = r22_out;
assign r4_write_en = 1'd1;
assign r4_clk = clk;
assign r4_reset = reset;
assign r4_in = r3_out;
assign r14_write_en = 1'd1;
assign r14_clk = clk;
assign r14_reset = reset;
assign r14_in = r13_out;
assign r2_write_en = 1'd1;
assign r2_clk = clk;
assign r2_reset = reset;
assign r2_in = r1_out;
assign r24_write_en = 1'd1;
assign r24_clk = clk;
assign r24_reset = reset;
assign r24_in = r23_out;
assign r17_write_en = 1'd1;
assign r17_clk = clk;
assign r17_reset = reset;
assign r17_in = r16_out;
assign r16_write_en = 1'd1;
assign r16_clk = clk;
assign r16_reset = reset;
assign r16_in = r15_out;
assign r3_write_en = 1'd1;
assign r3_clk = clk;
assign r3_reset = reset;
assign r3_in = r2_out;
assign r9_write_en = 1'd1;
assign r9_clk = clk;
assign r9_reset = reset;
assign r9_in = r8_out;
assign r21_write_en = 1'd1;
assign r21_clk = clk;
assign r21_reset = reset;
assign r21_in = r20_out;
assign r29_write_en = 1'd1;
assign r29_clk = clk;
assign r29_reset = reset;
assign r29_in = r28_out;
assign r6_write_en = 1'd1;
assign r6_clk = clk;
assign r6_reset = reset;
assign r6_in = r5_out;
assign r7_write_en = 1'd1;
assign r7_clk = clk;
assign r7_reset = reset;
assign r7_in = r6_out;
assign r8_write_en = 1'd1;
assign r8_clk = clk;
assign r8_reset = reset;
assign r8_in = r7_out;
// COMPONENT END: fsm_31
endmodule
module counter_128(
  input logic clk,
  input logic reset,
  output logic [6:0] state,
  output logic _0,
  input logic go,
  output logic done
);
// COMPONENT START: counter_128
logic [6:0] add_left;
logic [6:0] add_right;
logic [6:0] add_out;
logic [6:0] state0_in;
logic state0_write_en;
logic state0_clk;
logic state0_reset;
logic [6:0] state0_out;
logic state0_done;
logic done0_in;
logic done0_write_en;
logic done0_clk;
logic done0_reset;
logic done0_out;
logic done0_done;
std_add # (
    .WIDTH(7)
) add (
    .left(add_left),
    .out(add_out),
    .right(add_right)
);
std_reg # (
    .WIDTH(7)
) state0 (
    .clk(state0_clk),
    .done(state0_done),
    .in(state0_in),
    .out(state0_out),
    .reset(state0_reset),
    .write_en(state0_write_en)
);
std_reg # (
    .WIDTH(1)
) done0 (
    .clk(done0_clk),
    .done(done0_done),
    .in(done0_in),
    .out(done0_out),
    .reset(done0_reset),
    .write_en(done0_write_en)
);
wire _guard0 = 1;
wire _guard1 = go;
wire _guard2 = state0_out == 7'd0;
wire _guard3 = _guard1 & _guard2;
wire _guard4 = state0_out == 7'd127;
wire _guard5 = state0_out != 7'd127;
wire _guard6 = state0_out == 7'd127;
wire _guard7 = go;
wire _guard8 = state0_out != 7'd0;
wire _guard9 = _guard7 | _guard8;
wire _guard10 = state0_out != 7'd127;
wire _guard11 = _guard9 & _guard10;
wire _guard12 = _guard6 | _guard11;
wire _guard13 = state0_out == 7'd127;
wire _guard14 = go;
wire _guard15 = state0_out != 7'd0;
wire _guard16 = _guard14 | _guard15;
wire _guard17 = state0_out != 7'd127;
wire _guard18 = _guard16 & _guard17;
assign done = done0_out;
assign _0 = _guard3;
assign state = state0_out;
assign add_left = state0_out;
assign add_right = 7'd1;
assign done0_write_en = 1'd1;
assign done0_clk = clk;
assign done0_reset = reset;
assign done0_in =
  _guard4 ? 1'd1 :
  _guard5 ? 1'd0 :
  'x;
assign state0_write_en = _guard12;
assign state0_clk = clk;
assign state0_reset = reset;
assign state0_in =
  _guard13 ? 7'd0 :
  _guard18 ? add_out :
  'x;
// COMPONENT END: counter_128
endmodule
