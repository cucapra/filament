module ComplexMult_Exp8_Mant23(
  input wire clk,
  input wire [31:0] left_r,
  input wire [31:0] left_i,
  input wire [31:0] right_r,
  input wire [31:0] right_i,
  output wire [63:0] out
);
  // lint_off MULTIPLY
  function automatic [47:0] umul48b_24b_x_24b (input reg [23:0] lhs, input reg [23:0] rhs);
    begin
      umul48b_24b_x_24b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_left_r;
  reg [31:0] p0_left_i;
  reg [31:0] p0_right_r;
  reg [31:0] p0_right_i;
  always_ff @ (posedge clk) begin
    p0_left_r <= left_r;
    p0_left_i <= left_i;
    p0_right_r <= right_r;
    p0_right_i <= right_i;
  end

  // ===== Pipe stage 1:
  wire [22:0] p1_left_r_fraction__10_comb;
  wire [7:0] p1_left_r_bexp__9_comb;
  wire [22:0] p1_right_r_fraction__10_comb;
  wire [7:0] p1_right_r_bexp__9_comb;
  wire [22:0] p1_left_i_fraction__10_comb;
  wire [7:0] p1_left_i_bexp__9_comb;
  wire [22:0] p1_right_i_fraction__10_comb;
  wire [7:0] p1_right_i_bexp__9_comb;
  wire [23:0] p1_left_r_fraction__11_comb;
  wire [23:0] p1_right_r_fraction__11_comb;
  wire [23:0] p1_left_i_fraction__11_comb;
  wire [23:0] p1_right_i_fraction__11_comb;
  wire [8:0] p1_concat_4503_comb;
  wire [8:0] p1_concat_4504_comb;
  wire [23:0] p1_left_r_fraction__12_comb;
  wire [23:0] p1_right_r_fraction__12_comb;
  wire [8:0] p1_concat_4509_comb;
  wire [8:0] p1_concat_4510_comb;
  wire [23:0] p1_left_i_fraction__12_comb;
  wire [23:0] p1_right_i_fraction__12_comb;
  wire [8:0] p1_add_4516_comb;
  wire p1_eq_4517_comb;
  wire p1_eq_4518_comb;
  wire [47:0] p1_fraction__1_comb;
  wire [8:0] p1_add_4521_comb;
  wire p1_eq_4522_comb;
  wire p1_eq_4523_comb;
  wire [47:0] p1_fraction__8_comb;
  wire [8:0] p1_add_4526_comb;
  wire [47:0] p1_fraction__16_comb;
  wire [8:0] p1_add_4529_comb;
  wire [47:0] p1_fraction__24_comb;
  wire [9:0] p1_exp__1_comb;
  wire [47:0] p1_fraction__2_comb;
  wire [47:0] p1_sticky__1_comb;
  wire [9:0] p1_exp__4_comb;
  wire [47:0] p1_fraction__9_comb;
  wire [47:0] p1_sticky__2_comb;
  wire [9:0] p1_exp__8_comb;
  wire [47:0] p1_fraction__17_comb;
  wire [47:0] p1_sticky__4_comb;
  wire [9:0] p1_exp__12_comb;
  wire [47:0] p1_fraction__25_comb;
  wire [47:0] p1_sticky__6_comb;
  wire [9:0] p1_exp__2_comb;
  wire [47:0] p1_fraction__3_comb;
  wire [9:0] p1_exp__5_comb;
  wire [47:0] p1_fraction__10_comb;
  wire [9:0] p1_exp__9_comb;
  wire [47:0] p1_fraction__18_comb;
  wire [9:0] p1_exp__13_comb;
  wire [47:0] p1_fraction__26_comb;
  wire [9:0] p1_exp__3_comb;
  wire [9:0] p1_exp__6_comb;
  wire [9:0] p1_exp__10_comb;
  wire [9:0] p1_exp__14_comb;
  wire [47:0] p1_fraction__4_comb;
  wire [47:0] p1_sticky__5_comb;
  wire [47:0] p1_fraction__11_comb;
  wire [47:0] p1_sticky__3_comb;
  wire [47:0] p1_fraction__19_comb;
  wire [47:0] p1_sticky__7_comb;
  wire [47:0] p1_fraction__27_comb;
  wire [47:0] p1_sticky__8_comb;
  wire [47:0] p1_fraction__5_comb;
  wire [47:0] p1_fraction__12_comb;
  wire [47:0] p1_fraction__20_comb;
  wire [47:0] p1_fraction__28_comb;
  wire [7:0] p1_high_exp__6_comb;
  wire [7:0] p1_high_exp__1_comb;
  wire p1_eq_4735_comb;
  wire p1_eq_4737_comb;
  wire [7:0] p1_high_exp__3_comb;
  wire [7:0] p1_high_exp__4_comb;
  wire [22:0] p1_fraction__6_comb;
  wire [22:0] p1_fraction__13_comb;
  wire [22:0] p1_fraction__21_comb;
  wire [22:0] p1_fraction__29_comb;
  wire p1_and_4745_comb;
  wire p1_and_4746_comb;
  wire p1_eq_4731_comb;
  wire p1_eq_4733_comb;
  wire p1_greater_than_half_way__2_comb;
  wire [23:0] p1_fraction__7_comb;
  wire p1_greater_than_half_way__1_comb;
  wire [23:0] p1_fraction__14_comb;
  wire p1_greater_than_half_way__3_comb;
  wire [23:0] p1_fraction__22_comb;
  wire p1_greater_than_half_way__4_comb;
  wire [23:0] p1_fraction__30_comb;
  wire p1_has_0_arg__1_comb;
  wire p1_has_inf_arg__1_comb;
  wire p1_and_4741_comb;
  wire p1_and_4742_comb;
  wire p1_do_round_up__2_comb;
  wire [23:0] p1_add_4684_comb;
  wire p1_do_round_up__1_comb;
  wire [23:0] p1_add_4686_comb;
  wire p1_do_round_up__3_comb;
  wire [23:0] p1_add_4688_comb;
  wire p1_do_round_up__4_comb;
  wire [23:0] p1_add_4690_comb;
  wire p1_and_4764_comb;
  wire p1_and_4765_comb;
  wire p1_has_0_arg__2_comb;
  wire p1_has_inf_arg__2_comb;
  wire p1_has_0_arg__4_comb;
  wire p1_has_inf_arg__4_comb;
  wire p1_has_0_arg__3_comb;
  wire p1_has_inf_arg__3_comb;
  wire [23:0] p1_fraction__23_comb;
  wire [23:0] p1_fraction__15_comb;
  wire [23:0] p1_fraction__31_comb;
  wire [23:0] p1_fraction__32_comb;
  wire p1_is_result_nan__1_comb;
  wire p1_left_i_sign__2_comb;
  wire p1_right_i_sign__2_comb;
  wire p1_and_4760_comb;
  wire p1_and_4761_comb;
  wire [9:0] p1_add_4700_comb;
  wire [9:0] p1_add_4702_comb;
  wire [9:0] p1_add_4704_comb;
  wire [9:0] p1_add_4706_comb;
  wire p1_result_sign__2_comb;
  wire p1_is_result_nan__2_comb;
  wire p1_left_r_sign__2_comb;
  wire p1_right_r_sign__2_comb;
  wire p1_is_result_nan__4_comb;
  wire p1_is_result_nan__3_comb;
  wire [9:0] p1_exp__11_comb;
  wire [9:0] p1_exp__7_comb;
  wire [9:0] p1_exp__15_comb;
  wire [9:0] p1_exp__16_comb;
  wire p1_result_sign__3_comb;
  wire p1_result_sign__1_comb;
  wire p1_result_sign__6_comb;
  wire p1_result_sign__4_comb;
  wire p1_sgt_4715_comb;
  wire p1_sgt_4716_comb;
  wire p1_sgt_4717_comb;
  wire p1_sgt_4718_comb;
  wire [8:0] p1_result_exp__1_comb;
  wire [8:0] p1_result_exp__2_comb;
  wire [8:0] p1_result_exp__6_comb;
  wire [8:0] p1_result_exp__9_comb;
  wire p1_nor_4759_comb;
  wire p1_nor_4763_comb;
  wire p1_nor_4767_comb;
  wire p1_nor_4769_comb;
  wire [22:0] p1_result_fraction__3_comb;
  wire [22:0] p1_result_fraction__1_comb;
  wire [22:0] p1_result_fraction__6_comb;
  wire [22:0] p1_result_fraction__9_comb;
  wire p1_bd__1_sign_comb;
  wire p1_result_sign__5_comb;
  wire p1_result_sign__8_comb;
  wire p1_result_sign__7_comb;
  assign p1_left_r_fraction__10_comb = p0_left_r[22:0];
  assign p1_left_r_bexp__9_comb = p0_left_r[30:23];
  assign p1_right_r_fraction__10_comb = p0_right_r[22:0];
  assign p1_right_r_bexp__9_comb = p0_right_r[30:23];
  assign p1_left_i_fraction__10_comb = p0_left_i[22:0];
  assign p1_left_i_bexp__9_comb = p0_left_i[30:23];
  assign p1_right_i_fraction__10_comb = p0_right_i[22:0];
  assign p1_right_i_bexp__9_comb = p0_right_i[30:23];
  assign p1_left_r_fraction__11_comb = {1'h0, p1_left_r_fraction__10_comb} | 24'h80_0000;
  assign p1_right_r_fraction__11_comb = {1'h0, p1_right_r_fraction__10_comb} | 24'h80_0000;
  assign p1_left_i_fraction__11_comb = {1'h0, p1_left_i_fraction__10_comb} | 24'h80_0000;
  assign p1_right_i_fraction__11_comb = {1'h0, p1_right_i_fraction__10_comb} | 24'h80_0000;
  assign p1_concat_4503_comb = {1'h0, p1_left_r_bexp__9_comb};
  assign p1_concat_4504_comb = {1'h0, p1_right_r_bexp__9_comb};
  assign p1_left_r_fraction__12_comb = p1_left_r_fraction__11_comb & {24{p1_left_r_bexp__9_comb != 8'h00}};
  assign p1_right_r_fraction__12_comb = p1_right_r_fraction__11_comb & {24{p1_right_r_bexp__9_comb != 8'h00}};
  assign p1_concat_4509_comb = {1'h0, p1_left_i_bexp__9_comb};
  assign p1_concat_4510_comb = {1'h0, p1_right_i_bexp__9_comb};
  assign p1_left_i_fraction__12_comb = p1_left_i_fraction__11_comb & {24{p1_left_i_bexp__9_comb != 8'h00}};
  assign p1_right_i_fraction__12_comb = p1_right_i_fraction__11_comb & {24{p1_right_i_bexp__9_comb != 8'h00}};
  assign p1_add_4516_comb = p1_concat_4503_comb + p1_concat_4504_comb;
  assign p1_eq_4517_comb = p1_left_r_bexp__9_comb == 8'h00;
  assign p1_eq_4518_comb = p1_right_r_bexp__9_comb == 8'h00;
  assign p1_fraction__1_comb = umul48b_24b_x_24b(p1_left_r_fraction__12_comb, p1_right_r_fraction__12_comb);
  assign p1_add_4521_comb = p1_concat_4509_comb + p1_concat_4510_comb;
  assign p1_eq_4522_comb = p1_left_i_bexp__9_comb == 8'h00;
  assign p1_eq_4523_comb = p1_right_i_bexp__9_comb == 8'h00;
  assign p1_fraction__8_comb = umul48b_24b_x_24b(p1_left_i_fraction__12_comb, p1_right_i_fraction__12_comb);
  assign p1_add_4526_comb = p1_concat_4503_comb + p1_concat_4510_comb;
  assign p1_fraction__16_comb = umul48b_24b_x_24b(p1_left_r_fraction__12_comb, p1_right_i_fraction__12_comb);
  assign p1_add_4529_comb = p1_concat_4509_comb + p1_concat_4504_comb;
  assign p1_fraction__24_comb = umul48b_24b_x_24b(p1_left_i_fraction__12_comb, p1_right_r_fraction__12_comb);
  assign p1_exp__1_comb = {1'h0, p1_add_4516_comb} + 10'h381;
  assign p1_fraction__2_comb = p1_fraction__1_comb >> p1_fraction__1_comb[47];
  assign p1_sticky__1_comb = {47'h0000_0000_0000, p1_fraction__1_comb[0]};
  assign p1_exp__4_comb = {1'h0, p1_add_4521_comb} + 10'h381;
  assign p1_fraction__9_comb = p1_fraction__8_comb >> p1_fraction__8_comb[47];
  assign p1_sticky__2_comb = {47'h0000_0000_0000, p1_fraction__8_comb[0]};
  assign p1_exp__8_comb = {1'h0, p1_add_4526_comb} + 10'h381;
  assign p1_fraction__17_comb = p1_fraction__16_comb >> p1_fraction__16_comb[47];
  assign p1_sticky__4_comb = {47'h0000_0000_0000, p1_fraction__16_comb[0]};
  assign p1_exp__12_comb = {1'h0, p1_add_4529_comb} + 10'h381;
  assign p1_fraction__25_comb = p1_fraction__24_comb >> p1_fraction__24_comb[47];
  assign p1_sticky__6_comb = {47'h0000_0000_0000, p1_fraction__24_comb[0]};
  assign p1_exp__2_comb = p1_exp__1_comb & {10{~(p1_eq_4517_comb | p1_eq_4518_comb)}};
  assign p1_fraction__3_comb = p1_fraction__2_comb | p1_sticky__1_comb;
  assign p1_exp__5_comb = p1_exp__4_comb & {10{~(p1_eq_4522_comb | p1_eq_4523_comb)}};
  assign p1_fraction__10_comb = p1_fraction__9_comb | p1_sticky__2_comb;
  assign p1_exp__9_comb = p1_exp__8_comb & {10{~(p1_eq_4517_comb | p1_eq_4523_comb)}};
  assign p1_fraction__18_comb = p1_fraction__17_comb | p1_sticky__4_comb;
  assign p1_exp__13_comb = p1_exp__12_comb & {10{~(p1_eq_4522_comb | p1_eq_4518_comb)}};
  assign p1_fraction__26_comb = p1_fraction__25_comb | p1_sticky__6_comb;
  assign p1_exp__3_comb = p1_exp__2_comb + {9'h000, p1_fraction__1_comb[47]};
  assign p1_exp__6_comb = p1_exp__5_comb + {9'h000, p1_fraction__8_comb[47]};
  assign p1_exp__10_comb = p1_exp__9_comb + {9'h000, p1_fraction__16_comb[47]};
  assign p1_exp__14_comb = p1_exp__13_comb + {9'h000, p1_fraction__24_comb[47]};
  assign p1_fraction__4_comb = $signed(p1_exp__3_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__3_comb[47:1]} : p1_fraction__3_comb;
  assign p1_sticky__5_comb = {47'h0000_0000_0000, p1_fraction__3_comb[0]};
  assign p1_fraction__11_comb = $signed(p1_exp__6_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__10_comb[47:1]} : p1_fraction__10_comb;
  assign p1_sticky__3_comb = {47'h0000_0000_0000, p1_fraction__10_comb[0]};
  assign p1_fraction__19_comb = $signed(p1_exp__10_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__18_comb[47:1]} : p1_fraction__18_comb;
  assign p1_sticky__7_comb = {47'h0000_0000_0000, p1_fraction__18_comb[0]};
  assign p1_fraction__27_comb = $signed(p1_exp__14_comb) <= $signed(10'h000) ? {1'h0, p1_fraction__26_comb[47:1]} : p1_fraction__26_comb;
  assign p1_sticky__8_comb = {47'h0000_0000_0000, p1_fraction__26_comb[0]};
  assign p1_fraction__5_comb = p1_fraction__4_comb | p1_sticky__5_comb;
  assign p1_fraction__12_comb = p1_fraction__11_comb | p1_sticky__3_comb;
  assign p1_fraction__20_comb = p1_fraction__19_comb | p1_sticky__7_comb;
  assign p1_fraction__28_comb = p1_fraction__27_comb | p1_sticky__8_comb;
  assign p1_high_exp__6_comb = 8'hff;
  assign p1_high_exp__1_comb = 8'hff;
  assign p1_eq_4735_comb = p1_left_i_bexp__9_comb == p1_high_exp__6_comb;
  assign p1_eq_4737_comb = p1_right_i_bexp__9_comb == p1_high_exp__1_comb;
  assign p1_high_exp__3_comb = 8'hff;
  assign p1_high_exp__4_comb = 8'hff;
  assign p1_fraction__6_comb = p1_fraction__5_comb[45:23];
  assign p1_fraction__13_comb = p1_fraction__12_comb[45:23];
  assign p1_fraction__21_comb = p1_fraction__20_comb[45:23];
  assign p1_fraction__29_comb = p1_fraction__28_comb[45:23];
  assign p1_and_4745_comb = p1_eq_4735_comb & p1_left_i_fraction__10_comb == 23'h00_0000;
  assign p1_and_4746_comb = p1_eq_4737_comb & p1_right_i_fraction__10_comb == 23'h00_0000;
  assign p1_eq_4731_comb = p1_left_r_bexp__9_comb == p1_high_exp__3_comb;
  assign p1_eq_4733_comb = p1_right_r_bexp__9_comb == p1_high_exp__4_comb;
  assign p1_greater_than_half_way__2_comb = p1_fraction__5_comb[22] & p1_fraction__5_comb[21:0] != 22'h00_0000;
  assign p1_fraction__7_comb = {1'h0, p1_fraction__6_comb};
  assign p1_greater_than_half_way__1_comb = p1_fraction__12_comb[22] & p1_fraction__12_comb[21:0] != 22'h00_0000;
  assign p1_fraction__14_comb = {1'h0, p1_fraction__13_comb};
  assign p1_greater_than_half_way__3_comb = p1_fraction__20_comb[22] & p1_fraction__20_comb[21:0] != 22'h00_0000;
  assign p1_fraction__22_comb = {1'h0, p1_fraction__21_comb};
  assign p1_greater_than_half_way__4_comb = p1_fraction__28_comb[22] & p1_fraction__28_comb[21:0] != 22'h00_0000;
  assign p1_fraction__30_comb = {1'h0, p1_fraction__29_comb};
  assign p1_has_0_arg__1_comb = p1_eq_4522_comb | p1_eq_4523_comb;
  assign p1_has_inf_arg__1_comb = p1_and_4745_comb | p1_and_4746_comb;
  assign p1_and_4741_comb = p1_eq_4731_comb & p1_left_r_fraction__10_comb == 23'h00_0000;
  assign p1_and_4742_comb = p1_eq_4733_comb & p1_right_r_fraction__10_comb == 23'h00_0000;
  assign p1_do_round_up__2_comb = p1_greater_than_half_way__2_comb | p1_fraction__5_comb[22] & p1_fraction__5_comb[21:0] == 22'h00_0000 & p1_fraction__5_comb[23];
  assign p1_add_4684_comb = p1_fraction__7_comb + 24'h00_0001;
  assign p1_do_round_up__1_comb = p1_greater_than_half_way__1_comb | p1_fraction__12_comb[22] & p1_fraction__12_comb[21:0] == 22'h00_0000 & p1_fraction__12_comb[23];
  assign p1_add_4686_comb = p1_fraction__14_comb + 24'h00_0001;
  assign p1_do_round_up__3_comb = p1_greater_than_half_way__3_comb | p1_fraction__20_comb[22] & p1_fraction__20_comb[21:0] == 22'h00_0000 & p1_fraction__20_comb[23];
  assign p1_add_4688_comb = p1_fraction__22_comb + 24'h00_0001;
  assign p1_do_round_up__4_comb = p1_greater_than_half_way__4_comb | p1_fraction__28_comb[22] & p1_fraction__28_comb[21:0] == 22'h00_0000 & p1_fraction__28_comb[23];
  assign p1_add_4690_comb = p1_fraction__30_comb + 24'h00_0001;
  assign p1_and_4764_comb = p1_eq_4735_comb & p1_left_i_fraction__10_comb != 23'h00_0000;
  assign p1_and_4765_comb = p1_eq_4737_comb & p1_right_i_fraction__10_comb != 23'h00_0000;
  assign p1_has_0_arg__2_comb = p1_eq_4517_comb | p1_eq_4518_comb;
  assign p1_has_inf_arg__2_comb = p1_and_4741_comb | p1_and_4742_comb;
  assign p1_has_0_arg__4_comb = p1_eq_4522_comb | p1_eq_4518_comb;
  assign p1_has_inf_arg__4_comb = p1_and_4745_comb | p1_and_4742_comb;
  assign p1_has_0_arg__3_comb = p1_eq_4517_comb | p1_eq_4523_comb;
  assign p1_has_inf_arg__3_comb = p1_and_4741_comb | p1_and_4746_comb;
  assign p1_fraction__23_comb = p1_do_round_up__2_comb ? p1_add_4684_comb : p1_fraction__7_comb;
  assign p1_fraction__15_comb = p1_do_round_up__1_comb ? p1_add_4686_comb : p1_fraction__14_comb;
  assign p1_fraction__31_comb = p1_do_round_up__3_comb ? p1_add_4688_comb : p1_fraction__22_comb;
  assign p1_fraction__32_comb = p1_do_round_up__4_comb ? p1_add_4690_comb : p1_fraction__30_comb;
  assign p1_is_result_nan__1_comb = p1_and_4764_comb | p1_and_4765_comb | p1_has_0_arg__1_comb & p1_has_inf_arg__1_comb;
  assign p1_left_i_sign__2_comb = p0_left_i[31:31];
  assign p1_right_i_sign__2_comb = p0_right_i[31:31];
  assign p1_and_4760_comb = p1_eq_4731_comb & p1_left_r_fraction__10_comb != 23'h00_0000;
  assign p1_and_4761_comb = p1_eq_4733_comb & p1_right_r_fraction__10_comb != 23'h00_0000;
  assign p1_add_4700_comb = p1_exp__3_comb + 10'h001;
  assign p1_add_4702_comb = p1_exp__6_comb + 10'h001;
  assign p1_add_4704_comb = p1_exp__10_comb + 10'h001;
  assign p1_add_4706_comb = p1_exp__14_comb + 10'h001;
  assign p1_result_sign__2_comb = p1_left_i_sign__2_comb ^ p1_right_i_sign__2_comb;
  assign p1_is_result_nan__2_comb = p1_and_4760_comb | p1_and_4761_comb | p1_has_0_arg__2_comb & p1_has_inf_arg__2_comb;
  assign p1_left_r_sign__2_comb = p0_left_r[31:31];
  assign p1_right_r_sign__2_comb = p0_right_r[31:31];
  assign p1_is_result_nan__4_comb = p1_and_4764_comb | p1_and_4761_comb | p1_has_0_arg__4_comb & p1_has_inf_arg__4_comb;
  assign p1_is_result_nan__3_comb = p1_and_4760_comb | p1_and_4765_comb | p1_has_0_arg__3_comb & p1_has_inf_arg__3_comb;
  assign p1_exp__11_comb = p1_fraction__23_comb[23] ? p1_add_4700_comb : p1_exp__3_comb;
  assign p1_exp__7_comb = p1_fraction__15_comb[23] ? p1_add_4702_comb : p1_exp__6_comb;
  assign p1_exp__15_comb = p1_fraction__31_comb[23] ? p1_add_4704_comb : p1_exp__10_comb;
  assign p1_exp__16_comb = p1_fraction__32_comb[23] ? p1_add_4706_comb : p1_exp__14_comb;
  assign p1_result_sign__3_comb = ~p1_is_result_nan__1_comb & p1_result_sign__2_comb;
  assign p1_result_sign__1_comb = p1_left_r_sign__2_comb ^ p1_right_r_sign__2_comb;
  assign p1_result_sign__6_comb = p1_left_i_sign__2_comb ^ p1_right_r_sign__2_comb;
  assign p1_result_sign__4_comb = p1_left_r_sign__2_comb ^ p1_right_i_sign__2_comb;
  assign p1_sgt_4715_comb = $signed(p1_exp__11_comb) > $signed(10'h000);
  assign p1_sgt_4716_comb = $signed(p1_exp__7_comb) > $signed(10'h000);
  assign p1_sgt_4717_comb = $signed(p1_exp__15_comb) > $signed(10'h000);
  assign p1_sgt_4718_comb = $signed(p1_exp__16_comb) > $signed(10'h000);
  assign p1_result_exp__1_comb = p1_exp__11_comb[8:0];
  assign p1_result_exp__2_comb = p1_exp__7_comb[8:0];
  assign p1_result_exp__6_comb = p1_exp__15_comb[8:0];
  assign p1_result_exp__9_comb = p1_exp__16_comb[8:0];
  assign p1_nor_4759_comb = ~(p1_and_4741_comb | p1_and_4742_comb);
  assign p1_nor_4763_comb = ~(p1_and_4745_comb | p1_and_4746_comb);
  assign p1_nor_4767_comb = ~(p1_and_4741_comb | p1_and_4746_comb);
  assign p1_nor_4769_comb = ~(p1_and_4745_comb | p1_and_4742_comb);
  assign p1_result_fraction__3_comb = p1_fraction__23_comb[22:0];
  assign p1_result_fraction__1_comb = p1_fraction__15_comb[22:0];
  assign p1_result_fraction__6_comb = p1_fraction__31_comb[22:0];
  assign p1_result_fraction__9_comb = p1_fraction__32_comb[22:0];
  assign p1_bd__1_sign_comb = ~p1_result_sign__3_comb;
  assign p1_result_sign__5_comb = ~p1_is_result_nan__2_comb & p1_result_sign__1_comb;
  assign p1_result_sign__8_comb = ~p1_is_result_nan__4_comb & p1_result_sign__6_comb;
  assign p1_result_sign__7_comb = ~p1_is_result_nan__3_comb & p1_result_sign__4_comb;

  // Registers for pipe stage 1:
  reg p1_sgt_4715;
  reg p1_sgt_4716;
  reg p1_sgt_4717;
  reg p1_sgt_4718;
  reg [8:0] p1_result_exp__1;
  reg [8:0] p1_result_exp__2;
  reg [8:0] p1_result_exp__6;
  reg [8:0] p1_result_exp__9;
  reg p1_has_inf_arg__2;
  reg p1_has_inf_arg__1;
  reg p1_has_inf_arg__3;
  reg p1_has_inf_arg__4;
  reg p1_nor_4759;
  reg p1_nor_4763;
  reg p1_nor_4767;
  reg p1_nor_4769;
  reg [22:0] p1_result_fraction__3;
  reg p1_is_result_nan__2;
  reg [22:0] p1_result_fraction__1;
  reg p1_is_result_nan__1;
  reg [22:0] p1_result_fraction__6;
  reg p1_is_result_nan__3;
  reg [22:0] p1_result_fraction__9;
  reg p1_is_result_nan__4;
  reg p1_bd__1_sign;
  reg p1_result_sign__5;
  reg p1_result_sign__8;
  reg p1_result_sign__7;
  always_ff @ (posedge clk) begin
    p1_sgt_4715 <= p1_sgt_4715_comb;
    p1_sgt_4716 <= p1_sgt_4716_comb;
    p1_sgt_4717 <= p1_sgt_4717_comb;
    p1_sgt_4718 <= p1_sgt_4718_comb;
    p1_result_exp__1 <= p1_result_exp__1_comb;
    p1_result_exp__2 <= p1_result_exp__2_comb;
    p1_result_exp__6 <= p1_result_exp__6_comb;
    p1_result_exp__9 <= p1_result_exp__9_comb;
    p1_has_inf_arg__2 <= p1_has_inf_arg__2_comb;
    p1_has_inf_arg__1 <= p1_has_inf_arg__1_comb;
    p1_has_inf_arg__3 <= p1_has_inf_arg__3_comb;
    p1_has_inf_arg__4 <= p1_has_inf_arg__4_comb;
    p1_nor_4759 <= p1_nor_4759_comb;
    p1_nor_4763 <= p1_nor_4763_comb;
    p1_nor_4767 <= p1_nor_4767_comb;
    p1_nor_4769 <= p1_nor_4769_comb;
    p1_result_fraction__3 <= p1_result_fraction__3_comb;
    p1_is_result_nan__2 <= p1_is_result_nan__2_comb;
    p1_result_fraction__1 <= p1_result_fraction__1_comb;
    p1_is_result_nan__1 <= p1_is_result_nan__1_comb;
    p1_result_fraction__6 <= p1_result_fraction__6_comb;
    p1_is_result_nan__3 <= p1_is_result_nan__3_comb;
    p1_result_fraction__9 <= p1_result_fraction__9_comb;
    p1_is_result_nan__4 <= p1_is_result_nan__4_comb;
    p1_bd__1_sign <= p1_bd__1_sign_comb;
    p1_result_sign__5 <= p1_result_sign__5_comb;
    p1_result_sign__8 <= p1_result_sign__8_comb;
    p1_result_sign__7 <= p1_result_sign__7_comb;
  end

  // ===== Pipe stage 2:
  wire [8:0] p2_result_exp__4_comb;
  wire [8:0] p2_result_exp__3_comb;
  wire [8:0] p2_result_exp__7_comb;
  wire [8:0] p2_result_exp__10_comb;
  wire p2_nor_4903_comb;
  wire p2_nor_4904_comb;
  wire p2_nor_4905_comb;
  wire p2_nor_4906_comb;
  wire [22:0] p2_result_fraction__4_comb;
  wire [22:0] p2_nan_fraction__1_comb;
  wire [7:0] p2_high_exp__19_comb;
  wire [22:0] p2_result_fraction__2_comb;
  wire [22:0] p2_nan_fraction__5_comb;
  wire [7:0] p2_high_exp__18_comb;
  wire [22:0] p2_result_fraction__7_comb;
  wire [22:0] p2_nan_fraction__3_comb;
  wire [7:0] p2_high_exp__20_comb;
  wire [22:0] p2_result_fraction__10_comb;
  wire [22:0] p2_nan_fraction__4_comb;
  wire [7:0] p2_high_exp__21_comb;
  wire [22:0] p2_result_fraction__8_comb;
  wire [7:0] p2_result_exp__8_comb;
  wire [22:0] p2_result_fraction__5_comb;
  wire [7:0] p2_result_exp__5_comb;
  wire [22:0] p2_result_fraction__11_comb;
  wire [7:0] p2_result_exp__11_comb;
  wire [22:0] p2_result_fraction__12_comb;
  wire [7:0] p2_result_exp__12_comb;
  wire [5:0] p2_add_4978_comb;
  wire p2_ugt_4980_comb;
  wire [5:0] p2_add_4984_comb;
  wire [5:0] p2_add_4989_comb;
  wire p2_ugt_4991_comb;
  wire [5:0] p2_add_4995_comb;
  wire [27:0] p2_wide_x_comb;
  wire [7:0] p2_greater_exp_bexp_comb;
  wire [27:0] p2_wide_y_comb;
  wire [27:0] p2_wide_x__2_comb;
  wire [7:0] p2_greater_exp_bexp__1_comb;
  wire [27:0] p2_wide_y__2_comb;
  wire [27:0] p2_wide_x__1_comb;
  wire [7:0] p2_sub_5012_comb;
  wire [27:0] p2_wide_y__1_comb;
  wire [7:0] p2_sub_5014_comb;
  wire [27:0] p2_wide_x__3_comb;
  wire [7:0] p2_sub_5016_comb;
  wire [27:0] p2_wide_y__3_comb;
  wire [7:0] p2_sub_5018_comb;
  wire [27:0] p2_dropped_x_comb;
  wire [27:0] p2_dropped_y_comb;
  wire [27:0] p2_dropped_x__1_comb;
  wire [27:0] p2_dropped_y__1_comb;
  wire [7:0] p2_high_exp__22_comb;
  wire [7:0] p2_high_exp__23_comb;
  wire [7:0] p2_high_exp__24_comb;
  wire [7:0] p2_high_exp__25_comb;
  wire p2_eq_5077_comb;
  wire p2_eq_5078_comb;
  wire p2_eq_5079_comb;
  wire p2_eq_5080_comb;
  wire p2_eq_5081_comb;
  wire p2_eq_5082_comb;
  wire p2_eq_5083_comb;
  wire p2_eq_5084_comb;
  wire [7:0] p2_shift_x_comb;
  wire p2_sticky_x_comb;
  wire [7:0] p2_shift_y_comb;
  wire p2_sticky_y_comb;
  wire [7:0] p2_shift_x__1_comb;
  wire p2_sticky_x__1_comb;
  wire [7:0] p2_shift_y__1_comb;
  wire p2_sticky_y__1_comb;
  wire p2_and_5087_comb;
  wire p2_and_5088_comb;
  wire p2_and_5091_comb;
  wire p2_and_5092_comb;
  wire [27:0] p2_shifted_x_comb;
  wire [27:0] p2_shifted_y_comb;
  wire [27:0] p2_shifted_x__1_comb;
  wire [27:0] p2_shifted_y__1_comb;
  wire p2_greater_exp_sign_comb;
  wire [27:0] p2_addend_x_comb;
  wire [27:0] p2_addend_y_comb;
  wire p2_greater_exp_sign__1_comb;
  wire [27:0] p2_addend_x__2_comb;
  wire [27:0] p2_addend_y__2_comb;
  wire p2_has_pos_inf_comb;
  wire p2_has_neg_inf_comb;
  wire p2_has_pos_inf__1_comb;
  wire p2_has_neg_inf__1_comb;
  wire [27:0] p2_addend_x__1_comb;
  wire [27:0] p2_addend_y__1_comb;
  wire [27:0] p2_addend_x__3_comb;
  wire [27:0] p2_addend_y__3_comb;
  wire p2_nor_5116_comb;
  wire p2_nor_5120_comb;
  wire p2_is_result_nan__5_comb;
  wire p2_is_operand_inf_comb;
  wire p2_not_5123_comb;
  wire p2_is_result_nan__6_comb;
  wire p2_is_operand_inf__1_comb;
  wire p2_not_5126_comb;
  assign p2_result_exp__4_comb = p1_result_exp__1 & {9{p1_sgt_4715}};
  assign p2_result_exp__3_comb = p1_result_exp__2 & {9{p1_sgt_4716}};
  assign p2_result_exp__7_comb = p1_result_exp__6 & {9{p1_sgt_4717}};
  assign p2_result_exp__10_comb = p1_result_exp__9 & {9{p1_sgt_4718}};
  assign p2_nor_4903_comb = ~(p2_result_exp__4_comb[8] | p2_result_exp__4_comb[0] & p2_result_exp__4_comb[1] & p2_result_exp__4_comb[2] & p2_result_exp__4_comb[3] & p2_result_exp__4_comb[4] & p2_result_exp__4_comb[5] & p2_result_exp__4_comb[6] & p2_result_exp__4_comb[7]);
  assign p2_nor_4904_comb = ~(p2_result_exp__3_comb[8] | p2_result_exp__3_comb[0] & p2_result_exp__3_comb[1] & p2_result_exp__3_comb[2] & p2_result_exp__3_comb[3] & p2_result_exp__3_comb[4] & p2_result_exp__3_comb[5] & p2_result_exp__3_comb[6] & p2_result_exp__3_comb[7]);
  assign p2_nor_4905_comb = ~(p2_result_exp__7_comb[8] | p2_result_exp__7_comb[0] & p2_result_exp__7_comb[1] & p2_result_exp__7_comb[2] & p2_result_exp__7_comb[3] & p2_result_exp__7_comb[4] & p2_result_exp__7_comb[5] & p2_result_exp__7_comb[6] & p2_result_exp__7_comb[7]);
  assign p2_nor_4906_comb = ~(p2_result_exp__10_comb[8] | p2_result_exp__10_comb[0] & p2_result_exp__10_comb[1] & p2_result_exp__10_comb[2] & p2_result_exp__10_comb[3] & p2_result_exp__10_comb[4] & p2_result_exp__10_comb[5] & p2_result_exp__10_comb[6] & p2_result_exp__10_comb[7]);
  assign p2_result_fraction__4_comb = p1_result_fraction__3 & {23{p1_sgt_4715}} & {23{p2_nor_4903_comb}} & {23{p1_nor_4759}};
  assign p2_nan_fraction__1_comb = 23'h40_0000;
  assign p2_high_exp__19_comb = 8'hff;
  assign p2_result_fraction__2_comb = p1_result_fraction__1 & {23{p1_sgt_4716}} & {23{p2_nor_4904_comb}} & {23{p1_nor_4763}};
  assign p2_nan_fraction__5_comb = 23'h40_0000;
  assign p2_high_exp__18_comb = 8'hff;
  assign p2_result_fraction__7_comb = p1_result_fraction__6 & {23{p1_sgt_4717}} & {23{p2_nor_4905_comb}} & {23{p1_nor_4767}};
  assign p2_nan_fraction__3_comb = 23'h40_0000;
  assign p2_high_exp__20_comb = 8'hff;
  assign p2_result_fraction__10_comb = p1_result_fraction__9 & {23{p1_sgt_4718}} & {23{p2_nor_4906_comb}} & {23{p1_nor_4769}};
  assign p2_nan_fraction__4_comb = 23'h40_0000;
  assign p2_high_exp__21_comb = 8'hff;
  assign p2_result_fraction__8_comb = p1_is_result_nan__2 ? p2_nan_fraction__1_comb : p2_result_fraction__4_comb;
  assign p2_result_exp__8_comb = p1_is_result_nan__2 | p1_has_inf_arg__2 | ~p2_nor_4903_comb ? p2_high_exp__19_comb : p2_result_exp__4_comb[7:0];
  assign p2_result_fraction__5_comb = p1_is_result_nan__1 ? p2_nan_fraction__5_comb : p2_result_fraction__2_comb;
  assign p2_result_exp__5_comb = p1_is_result_nan__1 | p1_has_inf_arg__1 | ~p2_nor_4904_comb ? p2_high_exp__18_comb : p2_result_exp__3_comb[7:0];
  assign p2_result_fraction__11_comb = p1_is_result_nan__3 ? p2_nan_fraction__3_comb : p2_result_fraction__7_comb;
  assign p2_result_exp__11_comb = p1_is_result_nan__3 | p1_has_inf_arg__3 | ~p2_nor_4905_comb ? p2_high_exp__20_comb : p2_result_exp__7_comb[7:0];
  assign p2_result_fraction__12_comb = p1_is_result_nan__4 ? p2_nan_fraction__4_comb : p2_result_fraction__10_comb;
  assign p2_result_exp__12_comb = p1_is_result_nan__4 | p1_has_inf_arg__4 | ~p2_nor_4906_comb ? p2_high_exp__21_comb : p2_result_exp__10_comb[7:0];
  assign p2_add_4978_comb = p2_result_exp__8_comb[7:2] + 6'h07;
  assign p2_ugt_4980_comb = p2_result_exp__8_comb > p2_result_exp__5_comb;
  assign p2_add_4984_comb = p2_result_exp__5_comb[7:2] + 6'h07;
  assign p2_add_4989_comb = p2_result_exp__11_comb[7:2] + 6'h07;
  assign p2_ugt_4991_comb = p2_result_exp__11_comb > p2_result_exp__12_comb;
  assign p2_add_4995_comb = p2_result_exp__12_comb[7:2] + 6'h07;
  assign p2_wide_x_comb = {{2'h0, p2_result_fraction__8_comb} | 25'h080_0000, 3'h0};
  assign p2_greater_exp_bexp_comb = p2_ugt_4980_comb ? p2_result_exp__8_comb : p2_result_exp__5_comb;
  assign p2_wide_y_comb = {{2'h0, p2_result_fraction__5_comb} | 25'h080_0000, 3'h0};
  assign p2_wide_x__2_comb = {{2'h0, p2_result_fraction__11_comb} | 25'h080_0000, 3'h0};
  assign p2_greater_exp_bexp__1_comb = p2_ugt_4991_comb ? p2_result_exp__11_comb : p2_result_exp__12_comb;
  assign p2_wide_y__2_comb = {{2'h0, p2_result_fraction__12_comb} | 25'h080_0000, 3'h0};
  assign p2_wide_x__1_comb = p2_wide_x_comb & {28{p2_result_exp__8_comb != 8'h00}};
  assign p2_sub_5012_comb = {p2_add_4978_comb, p2_result_exp__8_comb[1:0]} - p2_greater_exp_bexp_comb;
  assign p2_wide_y__1_comb = p2_wide_y_comb & {28{p2_result_exp__5_comb != 8'h00}};
  assign p2_sub_5014_comb = {p2_add_4984_comb, p2_result_exp__5_comb[1:0]} - p2_greater_exp_bexp_comb;
  assign p2_wide_x__3_comb = p2_wide_x__2_comb & {28{p2_result_exp__11_comb != 8'h00}};
  assign p2_sub_5016_comb = {p2_add_4989_comb, p2_result_exp__11_comb[1:0]} - p2_greater_exp_bexp__1_comb;
  assign p2_wide_y__3_comb = p2_wide_y__2_comb & {28{p2_result_exp__12_comb != 8'h00}};
  assign p2_sub_5018_comb = {p2_add_4995_comb, p2_result_exp__12_comb[1:0]} - p2_greater_exp_bexp__1_comb;
  assign p2_dropped_x_comb = p2_sub_5012_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__1_comb << p2_sub_5012_comb;
  assign p2_dropped_y_comb = p2_sub_5014_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__1_comb << p2_sub_5014_comb;
  assign p2_dropped_x__1_comb = p2_sub_5016_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__3_comb << p2_sub_5016_comb;
  assign p2_dropped_y__1_comb = p2_sub_5018_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__3_comb << p2_sub_5018_comb;
  assign p2_high_exp__22_comb = 8'hff;
  assign p2_high_exp__23_comb = 8'hff;
  assign p2_high_exp__24_comb = 8'hff;
  assign p2_high_exp__25_comb = 8'hff;
  assign p2_eq_5077_comb = p2_result_exp__8_comb == p2_high_exp__22_comb;
  assign p2_eq_5078_comb = p2_result_fraction__8_comb == 23'h00_0000;
  assign p2_eq_5079_comb = p2_result_exp__5_comb == p2_high_exp__23_comb;
  assign p2_eq_5080_comb = p2_result_fraction__5_comb == 23'h00_0000;
  assign p2_eq_5081_comb = p2_result_exp__11_comb == p2_high_exp__24_comb;
  assign p2_eq_5082_comb = p2_result_fraction__11_comb == 23'h00_0000;
  assign p2_eq_5083_comb = p2_result_exp__12_comb == p2_high_exp__25_comb;
  assign p2_eq_5084_comb = p2_result_fraction__12_comb == 23'h00_0000;
  assign p2_shift_x_comb = p2_greater_exp_bexp_comb - p2_result_exp__8_comb;
  assign p2_sticky_x_comb = p2_dropped_x_comb[27:3] != 25'h000_0000;
  assign p2_shift_y_comb = p2_greater_exp_bexp_comb - p2_result_exp__5_comb;
  assign p2_sticky_y_comb = p2_dropped_y_comb[27:3] != 25'h000_0000;
  assign p2_shift_x__1_comb = p2_greater_exp_bexp__1_comb - p2_result_exp__11_comb;
  assign p2_sticky_x__1_comb = p2_dropped_x__1_comb[27:3] != 25'h000_0000;
  assign p2_shift_y__1_comb = p2_greater_exp_bexp__1_comb - p2_result_exp__12_comb;
  assign p2_sticky_y__1_comb = p2_dropped_y__1_comb[27:3] != 25'h000_0000;
  assign p2_and_5087_comb = p2_eq_5077_comb & p2_eq_5078_comb;
  assign p2_and_5088_comb = p2_eq_5079_comb & p2_eq_5080_comb;
  assign p2_and_5091_comb = p2_eq_5081_comb & p2_eq_5082_comb;
  assign p2_and_5092_comb = p2_eq_5083_comb & p2_eq_5084_comb;
  assign p2_shifted_x_comb = p2_shift_x_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__1_comb >> p2_shift_x_comb;
  assign p2_shifted_y_comb = p2_shift_y_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__1_comb >> p2_shift_y_comb;
  assign p2_shifted_x__1_comb = p2_shift_x__1_comb >= 8'h1c ? 28'h000_0000 : p2_wide_x__3_comb >> p2_shift_x__1_comb;
  assign p2_shifted_y__1_comb = p2_shift_y__1_comb >= 8'h1c ? 28'h000_0000 : p2_wide_y__3_comb >> p2_shift_y__1_comb;
  assign p2_greater_exp_sign_comb = p2_ugt_4980_comb ? p1_result_sign__5 : p1_bd__1_sign;
  assign p2_addend_x_comb = p2_shifted_x_comb | {27'h000_0000, p2_sticky_x_comb};
  assign p2_addend_y_comb = p2_shifted_y_comb | {27'h000_0000, p2_sticky_y_comb};
  assign p2_greater_exp_sign__1_comb = p2_ugt_4991_comb ? p1_result_sign__7 : p1_result_sign__8;
  assign p2_addend_x__2_comb = p2_shifted_x__1_comb | {27'h000_0000, p2_sticky_x__1_comb};
  assign p2_addend_y__2_comb = p2_shifted_y__1_comb | {27'h000_0000, p2_sticky_y__1_comb};
  assign p2_has_pos_inf_comb = ~(~(p2_eq_5077_comb & p2_eq_5078_comb) | p1_result_sign__5) | ~(~(p2_eq_5079_comb & p2_eq_5080_comb) | p1_bd__1_sign);
  assign p2_has_neg_inf_comb = p2_and_5087_comb & p1_result_sign__5 | p2_and_5088_comb & p1_bd__1_sign;
  assign p2_has_pos_inf__1_comb = ~(~(p2_eq_5081_comb & p2_eq_5082_comb) | p1_result_sign__7) | ~(~(p2_eq_5083_comb & p2_eq_5084_comb) | p1_result_sign__8);
  assign p2_has_neg_inf__1_comb = p2_and_5091_comb & p1_result_sign__7 | p2_and_5092_comb & p1_result_sign__8;
  assign p2_addend_x__1_comb = p1_result_sign__5 ^ p2_greater_exp_sign_comb ? -p2_addend_x_comb : p2_addend_x_comb;
  assign p2_addend_y__1_comb = p1_bd__1_sign ^ p2_greater_exp_sign_comb ? -p2_addend_y_comb : p2_addend_y_comb;
  assign p2_addend_x__3_comb = p1_result_sign__7 ^ p2_greater_exp_sign__1_comb ? -p2_addend_x__2_comb : p2_addend_x__2_comb;
  assign p2_addend_y__3_comb = p1_result_sign__8 ^ p2_greater_exp_sign__1_comb ? -p2_addend_y__2_comb : p2_addend_y__2_comb;
  assign p2_nor_5116_comb = ~(p2_and_5087_comb | p2_and_5088_comb);
  assign p2_nor_5120_comb = ~(p2_and_5091_comb | p2_and_5092_comb);
  assign p2_is_result_nan__5_comb = p2_eq_5077_comb & p2_result_fraction__8_comb != 23'h00_0000 | p2_eq_5079_comb & p2_result_fraction__5_comb != 23'h00_0000 | p2_has_pos_inf_comb & p2_has_neg_inf_comb;
  assign p2_is_operand_inf_comb = p2_and_5087_comb | p2_and_5088_comb;
  assign p2_not_5123_comb = ~p2_has_pos_inf_comb;
  assign p2_is_result_nan__6_comb = p2_eq_5081_comb & p2_result_fraction__11_comb != 23'h00_0000 | p2_eq_5083_comb & p2_result_fraction__12_comb != 23'h00_0000 | p2_has_pos_inf__1_comb & p2_has_neg_inf__1_comb;
  assign p2_is_operand_inf__1_comb = p2_and_5091_comb | p2_and_5092_comb;
  assign p2_not_5126_comb = ~p2_has_pos_inf__1_comb;

  // Registers for pipe stage 2:
  reg [7:0] p2_greater_exp_bexp;
  reg [7:0] p2_greater_exp_bexp__1;
  reg p2_greater_exp_sign;
  reg p2_greater_exp_sign__1;
  reg [27:0] p2_addend_x__1;
  reg [27:0] p2_addend_y__1;
  reg [27:0] p2_addend_x__3;
  reg [27:0] p2_addend_y__3;
  reg p2_nor_5116;
  reg p2_nor_5120;
  reg p2_is_result_nan__5;
  reg p2_is_operand_inf;
  reg p2_not_5123;
  reg p2_is_result_nan__6;
  reg p2_is_operand_inf__1;
  reg p2_not_5126;
  always_ff @ (posedge clk) begin
    p2_greater_exp_bexp <= p2_greater_exp_bexp_comb;
    p2_greater_exp_bexp__1 <= p2_greater_exp_bexp__1_comb;
    p2_greater_exp_sign <= p2_greater_exp_sign_comb;
    p2_greater_exp_sign__1 <= p2_greater_exp_sign__1_comb;
    p2_addend_x__1 <= p2_addend_x__1_comb;
    p2_addend_y__1 <= p2_addend_y__1_comb;
    p2_addend_x__3 <= p2_addend_x__3_comb;
    p2_addend_y__3 <= p2_addend_y__3_comb;
    p2_nor_5116 <= p2_nor_5116_comb;
    p2_nor_5120 <= p2_nor_5120_comb;
    p2_is_result_nan__5 <= p2_is_result_nan__5_comb;
    p2_is_operand_inf <= p2_is_operand_inf_comb;
    p2_not_5123 <= p2_not_5123_comb;
    p2_is_result_nan__6 <= p2_is_result_nan__6_comb;
    p2_is_operand_inf__1 <= p2_is_operand_inf__1_comb;
    p2_not_5126 <= p2_not_5126_comb;
  end

  // ===== Pipe stage 3:
  wire [28:0] p3_fraction__33_comb;
  wire [28:0] p3_fraction__34_comb;
  wire [27:0] p3_abs_fraction_comb;
  wire [27:0] p3_abs_fraction__1_comb;
  wire [27:0] p3_reverse_5175_comb;
  wire [27:0] p3_reverse_5176_comb;
  wire [28:0] p3_one_hot_5177_comb;
  wire [28:0] p3_one_hot_5178_comb;
  wire [4:0] p3_encode_5179_comb;
  wire [4:0] p3_encode_5180_comb;
  wire p3_carry_bit_comb;
  wire p3_cancel_comb;
  wire p3_carry_bit__1_comb;
  wire p3_cancel__1_comb;
  wire [27:0] p3_leading_zeroes_comb;
  wire [27:0] p3_leading_zeroes__1_comb;
  wire p3_and_5207_comb;
  wire p3_and_5208_comb;
  wire p3_and_5209_comb;
  wire [26:0] p3_carry_fraction_comb;
  wire [27:0] p3_add_5213_comb;
  wire p3_and_5214_comb;
  wire p3_and_5215_comb;
  wire p3_and_5216_comb;
  wire [26:0] p3_carry_fraction__2_comb;
  wire [27:0] p3_add_5220_comb;
  wire [2:0] p3_concat_5221_comb;
  wire [26:0] p3_carry_fraction__1_comb;
  wire [26:0] p3_cancel_fraction_comb;
  wire [2:0] p3_concat_5224_comb;
  wire [26:0] p3_carry_fraction__3_comb;
  wire [26:0] p3_cancel_fraction__1_comb;
  wire [26:0] p3_shifted_fraction_comb;
  wire [26:0] p3_shifted_fraction__1_comb;
  wire p3_fraction_is_zero_comb;
  wire p3_fraction_is_zero__1_comb;
  wire [2:0] p3_normal_chunk_comb;
  wire [1:0] p3_half_way_chunk_comb;
  wire [2:0] p3_normal_chunk__1_comb;
  wire [1:0] p3_half_way_chunk__1_comb;
  wire [24:0] p3_add_5248_comb;
  wire [24:0] p3_add_5252_comb;
  wire p3_result_sign__9_comb;
  wire p3_result_sign__11_comb;
  wire p3_do_round_up__5_comb;
  wire p3_do_round_up__6_comb;
  wire p3_result_sign__10_comb;
  wire p3_result_sign__12_comb;
  wire [27:0] p3_rounded_fraction_comb;
  wire [27:0] p3_rounded_fraction__1_comb;
  wire p3_ne_5263_comb;
  wire p3_ne_5264_comb;
  wire p3_result_sign__13_comb;
  wire p3_result_sign__14_comb;
  assign p3_fraction__33_comb = {{1{p2_addend_x__1[27]}}, p2_addend_x__1} + {{1{p2_addend_y__1[27]}}, p2_addend_y__1};
  assign p3_fraction__34_comb = {{1{p2_addend_x__3[27]}}, p2_addend_x__3} + {{1{p2_addend_y__3[27]}}, p2_addend_y__3};
  assign p3_abs_fraction_comb = p3_fraction__33_comb[28] ? -p3_fraction__33_comb[27:0] : p3_fraction__33_comb[27:0];
  assign p3_abs_fraction__1_comb = p3_fraction__34_comb[28] ? -p3_fraction__34_comb[27:0] : p3_fraction__34_comb[27:0];
  assign p3_reverse_5175_comb = {p3_abs_fraction_comb[0], p3_abs_fraction_comb[1], p3_abs_fraction_comb[2], p3_abs_fraction_comb[3], p3_abs_fraction_comb[4], p3_abs_fraction_comb[5], p3_abs_fraction_comb[6], p3_abs_fraction_comb[7], p3_abs_fraction_comb[8], p3_abs_fraction_comb[9], p3_abs_fraction_comb[10], p3_abs_fraction_comb[11], p3_abs_fraction_comb[12], p3_abs_fraction_comb[13], p3_abs_fraction_comb[14], p3_abs_fraction_comb[15], p3_abs_fraction_comb[16], p3_abs_fraction_comb[17], p3_abs_fraction_comb[18], p3_abs_fraction_comb[19], p3_abs_fraction_comb[20], p3_abs_fraction_comb[21], p3_abs_fraction_comb[22], p3_abs_fraction_comb[23], p3_abs_fraction_comb[24], p3_abs_fraction_comb[25], p3_abs_fraction_comb[26], p3_abs_fraction_comb[27]};
  assign p3_reverse_5176_comb = {p3_abs_fraction__1_comb[0], p3_abs_fraction__1_comb[1], p3_abs_fraction__1_comb[2], p3_abs_fraction__1_comb[3], p3_abs_fraction__1_comb[4], p3_abs_fraction__1_comb[5], p3_abs_fraction__1_comb[6], p3_abs_fraction__1_comb[7], p3_abs_fraction__1_comb[8], p3_abs_fraction__1_comb[9], p3_abs_fraction__1_comb[10], p3_abs_fraction__1_comb[11], p3_abs_fraction__1_comb[12], p3_abs_fraction__1_comb[13], p3_abs_fraction__1_comb[14], p3_abs_fraction__1_comb[15], p3_abs_fraction__1_comb[16], p3_abs_fraction__1_comb[17], p3_abs_fraction__1_comb[18], p3_abs_fraction__1_comb[19], p3_abs_fraction__1_comb[20], p3_abs_fraction__1_comb[21], p3_abs_fraction__1_comb[22], p3_abs_fraction__1_comb[23], p3_abs_fraction__1_comb[24], p3_abs_fraction__1_comb[25], p3_abs_fraction__1_comb[26], p3_abs_fraction__1_comb[27]};
  assign p3_one_hot_5177_comb = {p3_reverse_5175_comb[27:0] == 28'h000_0000, p3_reverse_5175_comb[27] && p3_reverse_5175_comb[26:0] == 27'h000_0000, p3_reverse_5175_comb[26] && p3_reverse_5175_comb[25:0] == 26'h000_0000, p3_reverse_5175_comb[25] && p3_reverse_5175_comb[24:0] == 25'h000_0000, p3_reverse_5175_comb[24] && p3_reverse_5175_comb[23:0] == 24'h00_0000, p3_reverse_5175_comb[23] && p3_reverse_5175_comb[22:0] == 23'h00_0000, p3_reverse_5175_comb[22] && p3_reverse_5175_comb[21:0] == 22'h00_0000, p3_reverse_5175_comb[21] && p3_reverse_5175_comb[20:0] == 21'h00_0000, p3_reverse_5175_comb[20] && p3_reverse_5175_comb[19:0] == 20'h0_0000, p3_reverse_5175_comb[19] && p3_reverse_5175_comb[18:0] == 19'h0_0000, p3_reverse_5175_comb[18] && p3_reverse_5175_comb[17:0] == 18'h0_0000, p3_reverse_5175_comb[17] && p3_reverse_5175_comb[16:0] == 17'h0_0000, p3_reverse_5175_comb[16] && p3_reverse_5175_comb[15:0] == 16'h0000, p3_reverse_5175_comb[15] && p3_reverse_5175_comb[14:0] == 15'h0000, p3_reverse_5175_comb[14] && p3_reverse_5175_comb[13:0] == 14'h0000, p3_reverse_5175_comb[13] && p3_reverse_5175_comb[12:0] == 13'h0000, p3_reverse_5175_comb[12] && p3_reverse_5175_comb[11:0] == 12'h000, p3_reverse_5175_comb[11] && p3_reverse_5175_comb[10:0] == 11'h000, p3_reverse_5175_comb[10] && p3_reverse_5175_comb[9:0] == 10'h000, p3_reverse_5175_comb[9] && p3_reverse_5175_comb[8:0] == 9'h000, p3_reverse_5175_comb[8] && p3_reverse_5175_comb[7:0] == 8'h00, p3_reverse_5175_comb[7] && p3_reverse_5175_comb[6:0] == 7'h00, p3_reverse_5175_comb[6] && p3_reverse_5175_comb[5:0] == 6'h00, p3_reverse_5175_comb[5] && p3_reverse_5175_comb[4:0] == 5'h00, p3_reverse_5175_comb[4] && p3_reverse_5175_comb[3:0] == 4'h0, p3_reverse_5175_comb[3] && p3_reverse_5175_comb[2:0] == 3'h0, p3_reverse_5175_comb[2] && p3_reverse_5175_comb[1:0] == 2'h0, p3_reverse_5175_comb[1] && !p3_reverse_5175_comb[0], p3_reverse_5175_comb[0]};
  assign p3_one_hot_5178_comb = {p3_reverse_5176_comb[27:0] == 28'h000_0000, p3_reverse_5176_comb[27] && p3_reverse_5176_comb[26:0] == 27'h000_0000, p3_reverse_5176_comb[26] && p3_reverse_5176_comb[25:0] == 26'h000_0000, p3_reverse_5176_comb[25] && p3_reverse_5176_comb[24:0] == 25'h000_0000, p3_reverse_5176_comb[24] && p3_reverse_5176_comb[23:0] == 24'h00_0000, p3_reverse_5176_comb[23] && p3_reverse_5176_comb[22:0] == 23'h00_0000, p3_reverse_5176_comb[22] && p3_reverse_5176_comb[21:0] == 22'h00_0000, p3_reverse_5176_comb[21] && p3_reverse_5176_comb[20:0] == 21'h00_0000, p3_reverse_5176_comb[20] && p3_reverse_5176_comb[19:0] == 20'h0_0000, p3_reverse_5176_comb[19] && p3_reverse_5176_comb[18:0] == 19'h0_0000, p3_reverse_5176_comb[18] && p3_reverse_5176_comb[17:0] == 18'h0_0000, p3_reverse_5176_comb[17] && p3_reverse_5176_comb[16:0] == 17'h0_0000, p3_reverse_5176_comb[16] && p3_reverse_5176_comb[15:0] == 16'h0000, p3_reverse_5176_comb[15] && p3_reverse_5176_comb[14:0] == 15'h0000, p3_reverse_5176_comb[14] && p3_reverse_5176_comb[13:0] == 14'h0000, p3_reverse_5176_comb[13] && p3_reverse_5176_comb[12:0] == 13'h0000, p3_reverse_5176_comb[12] && p3_reverse_5176_comb[11:0] == 12'h000, p3_reverse_5176_comb[11] && p3_reverse_5176_comb[10:0] == 11'h000, p3_reverse_5176_comb[10] && p3_reverse_5176_comb[9:0] == 10'h000, p3_reverse_5176_comb[9] && p3_reverse_5176_comb[8:0] == 9'h000, p3_reverse_5176_comb[8] && p3_reverse_5176_comb[7:0] == 8'h00, p3_reverse_5176_comb[7] && p3_reverse_5176_comb[6:0] == 7'h00, p3_reverse_5176_comb[6] && p3_reverse_5176_comb[5:0] == 6'h00, p3_reverse_5176_comb[5] && p3_reverse_5176_comb[4:0] == 5'h00, p3_reverse_5176_comb[4] && p3_reverse_5176_comb[3:0] == 4'h0, p3_reverse_5176_comb[3] && p3_reverse_5176_comb[2:0] == 3'h0, p3_reverse_5176_comb[2] && p3_reverse_5176_comb[1:0] == 2'h0, p3_reverse_5176_comb[1] && !p3_reverse_5176_comb[0], p3_reverse_5176_comb[0]};
  assign p3_encode_5179_comb = {p3_one_hot_5177_comb[16] | p3_one_hot_5177_comb[17] | p3_one_hot_5177_comb[18] | p3_one_hot_5177_comb[19] | p3_one_hot_5177_comb[20] | p3_one_hot_5177_comb[21] | p3_one_hot_5177_comb[22] | p3_one_hot_5177_comb[23] | p3_one_hot_5177_comb[24] | p3_one_hot_5177_comb[25] | p3_one_hot_5177_comb[26] | p3_one_hot_5177_comb[27] | p3_one_hot_5177_comb[28], p3_one_hot_5177_comb[8] | p3_one_hot_5177_comb[9] | p3_one_hot_5177_comb[10] | p3_one_hot_5177_comb[11] | p3_one_hot_5177_comb[12] | p3_one_hot_5177_comb[13] | p3_one_hot_5177_comb[14] | p3_one_hot_5177_comb[15] | p3_one_hot_5177_comb[24] | p3_one_hot_5177_comb[25] | p3_one_hot_5177_comb[26] | p3_one_hot_5177_comb[27] | p3_one_hot_5177_comb[28], p3_one_hot_5177_comb[4] | p3_one_hot_5177_comb[5] | p3_one_hot_5177_comb[6] | p3_one_hot_5177_comb[7] | p3_one_hot_5177_comb[12] | p3_one_hot_5177_comb[13] | p3_one_hot_5177_comb[14] | p3_one_hot_5177_comb[15] | p3_one_hot_5177_comb[20] | p3_one_hot_5177_comb[21] | p3_one_hot_5177_comb[22] | p3_one_hot_5177_comb[23] | p3_one_hot_5177_comb[28], p3_one_hot_5177_comb[2] | p3_one_hot_5177_comb[3] | p3_one_hot_5177_comb[6] | p3_one_hot_5177_comb[7] | p3_one_hot_5177_comb[10] | p3_one_hot_5177_comb[11] | p3_one_hot_5177_comb[14] | p3_one_hot_5177_comb[15] | p3_one_hot_5177_comb[18] | p3_one_hot_5177_comb[19] | p3_one_hot_5177_comb[22] | p3_one_hot_5177_comb[23] | p3_one_hot_5177_comb[26] | p3_one_hot_5177_comb[27], p3_one_hot_5177_comb[1] | p3_one_hot_5177_comb[3] | p3_one_hot_5177_comb[5] | p3_one_hot_5177_comb[7] | p3_one_hot_5177_comb[9] | p3_one_hot_5177_comb[11] | p3_one_hot_5177_comb[13] | p3_one_hot_5177_comb[15] | p3_one_hot_5177_comb[17] | p3_one_hot_5177_comb[19] | p3_one_hot_5177_comb[21] | p3_one_hot_5177_comb[23] | p3_one_hot_5177_comb[25] | p3_one_hot_5177_comb[27]};
  assign p3_encode_5180_comb = {p3_one_hot_5178_comb[16] | p3_one_hot_5178_comb[17] | p3_one_hot_5178_comb[18] | p3_one_hot_5178_comb[19] | p3_one_hot_5178_comb[20] | p3_one_hot_5178_comb[21] | p3_one_hot_5178_comb[22] | p3_one_hot_5178_comb[23] | p3_one_hot_5178_comb[24] | p3_one_hot_5178_comb[25] | p3_one_hot_5178_comb[26] | p3_one_hot_5178_comb[27] | p3_one_hot_5178_comb[28], p3_one_hot_5178_comb[8] | p3_one_hot_5178_comb[9] | p3_one_hot_5178_comb[10] | p3_one_hot_5178_comb[11] | p3_one_hot_5178_comb[12] | p3_one_hot_5178_comb[13] | p3_one_hot_5178_comb[14] | p3_one_hot_5178_comb[15] | p3_one_hot_5178_comb[24] | p3_one_hot_5178_comb[25] | p3_one_hot_5178_comb[26] | p3_one_hot_5178_comb[27] | p3_one_hot_5178_comb[28], p3_one_hot_5178_comb[4] | p3_one_hot_5178_comb[5] | p3_one_hot_5178_comb[6] | p3_one_hot_5178_comb[7] | p3_one_hot_5178_comb[12] | p3_one_hot_5178_comb[13] | p3_one_hot_5178_comb[14] | p3_one_hot_5178_comb[15] | p3_one_hot_5178_comb[20] | p3_one_hot_5178_comb[21] | p3_one_hot_5178_comb[22] | p3_one_hot_5178_comb[23] | p3_one_hot_5178_comb[28], p3_one_hot_5178_comb[2] | p3_one_hot_5178_comb[3] | p3_one_hot_5178_comb[6] | p3_one_hot_5178_comb[7] | p3_one_hot_5178_comb[10] | p3_one_hot_5178_comb[11] | p3_one_hot_5178_comb[14] | p3_one_hot_5178_comb[15] | p3_one_hot_5178_comb[18] | p3_one_hot_5178_comb[19] | p3_one_hot_5178_comb[22] | p3_one_hot_5178_comb[23] | p3_one_hot_5178_comb[26] | p3_one_hot_5178_comb[27], p3_one_hot_5178_comb[1] | p3_one_hot_5178_comb[3] | p3_one_hot_5178_comb[5] | p3_one_hot_5178_comb[7] | p3_one_hot_5178_comb[9] | p3_one_hot_5178_comb[11] | p3_one_hot_5178_comb[13] | p3_one_hot_5178_comb[15] | p3_one_hot_5178_comb[17] | p3_one_hot_5178_comb[19] | p3_one_hot_5178_comb[21] | p3_one_hot_5178_comb[23] | p3_one_hot_5178_comb[25] | p3_one_hot_5178_comb[27]};
  assign p3_carry_bit_comb = p3_abs_fraction_comb[27];
  assign p3_cancel_comb = p3_encode_5179_comb[1] | p3_encode_5179_comb[2] | p3_encode_5179_comb[3] | p3_encode_5179_comb[4];
  assign p3_carry_bit__1_comb = p3_abs_fraction__1_comb[27];
  assign p3_cancel__1_comb = p3_encode_5180_comb[1] | p3_encode_5180_comb[2] | p3_encode_5180_comb[3] | p3_encode_5180_comb[4];
  assign p3_leading_zeroes_comb = {23'h00_0000, p3_encode_5179_comb};
  assign p3_leading_zeroes__1_comb = {23'h00_0000, p3_encode_5180_comb};
  assign p3_and_5207_comb = ~p3_carry_bit_comb & ~p3_cancel_comb;
  assign p3_and_5208_comb = ~p3_carry_bit_comb & p3_cancel_comb;
  assign p3_and_5209_comb = p3_carry_bit_comb & ~p3_cancel_comb;
  assign p3_carry_fraction_comb = p3_abs_fraction_comb[27:1];
  assign p3_add_5213_comb = p3_leading_zeroes_comb + 28'hfff_ffff;
  assign p3_and_5214_comb = ~p3_carry_bit__1_comb & ~p3_cancel__1_comb;
  assign p3_and_5215_comb = ~p3_carry_bit__1_comb & p3_cancel__1_comb;
  assign p3_and_5216_comb = p3_carry_bit__1_comb & ~p3_cancel__1_comb;
  assign p3_carry_fraction__2_comb = p3_abs_fraction__1_comb[27:1];
  assign p3_add_5220_comb = p3_leading_zeroes__1_comb + 28'hfff_ffff;
  assign p3_concat_5221_comb = {p3_and_5207_comb, p3_and_5208_comb, p3_and_5209_comb};
  assign p3_carry_fraction__1_comb = p3_carry_fraction_comb | {26'h000_0000, p3_abs_fraction_comb[0]};
  assign p3_cancel_fraction_comb = p3_add_5213_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction_comb[26:0] << p3_add_5213_comb;
  assign p3_concat_5224_comb = {p3_and_5214_comb, p3_and_5215_comb, p3_and_5216_comb};
  assign p3_carry_fraction__3_comb = p3_carry_fraction__2_comb | {26'h000_0000, p3_abs_fraction__1_comb[0]};
  assign p3_cancel_fraction__1_comb = p3_add_5220_comb >= 28'h000_001b ? 27'h000_0000 : p3_abs_fraction__1_comb[26:0] << p3_add_5220_comb;
  assign p3_shifted_fraction_comb = p3_carry_fraction__1_comb & {27{p3_concat_5221_comb[0]}} | p3_cancel_fraction_comb & {27{p3_concat_5221_comb[1]}} | p3_abs_fraction_comb[26:0] & {27{p3_concat_5221_comb[2]}};
  assign p3_shifted_fraction__1_comb = p3_carry_fraction__3_comb & {27{p3_concat_5224_comb[0]}} | p3_cancel_fraction__1_comb & {27{p3_concat_5224_comb[1]}} | p3_abs_fraction__1_comb[26:0] & {27{p3_concat_5224_comb[2]}};
  assign p3_fraction_is_zero_comb = p3_fraction__33_comb == 29'h0000_0000;
  assign p3_fraction_is_zero__1_comb = p3_fraction__34_comb == 29'h0000_0000;
  assign p3_normal_chunk_comb = p3_shifted_fraction_comb[2:0];
  assign p3_half_way_chunk_comb = p3_shifted_fraction_comb[3:2];
  assign p3_normal_chunk__1_comb = p3_shifted_fraction__1_comb[2:0];
  assign p3_half_way_chunk__1_comb = p3_shifted_fraction__1_comb[3:2];
  assign p3_add_5248_comb = {1'h0, p3_shifted_fraction_comb[26:3]} + 25'h000_0001;
  assign p3_add_5252_comb = {1'h0, p3_shifted_fraction__1_comb[26:3]} + 25'h000_0001;
  assign p3_result_sign__9_comb = ~(~p3_fraction__33_comb[28] | p2_greater_exp_sign) | ~(p3_fraction__33_comb[28] | p3_fraction_is_zero_comb | ~p2_greater_exp_sign);
  assign p3_result_sign__11_comb = ~(~p3_fraction__34_comb[28] | p2_greater_exp_sign__1) | ~(p3_fraction__34_comb[28] | p3_fraction_is_zero__1_comb | ~p2_greater_exp_sign__1);
  assign p3_do_round_up__5_comb = p3_normal_chunk_comb > 3'h4 | p3_half_way_chunk_comb == 2'h3;
  assign p3_do_round_up__6_comb = p3_normal_chunk__1_comb > 3'h4 | p3_half_way_chunk__1_comb == 2'h3;
  assign p3_result_sign__10_comb = p2_is_operand_inf ? p2_not_5123 : p3_result_sign__9_comb;
  assign p3_result_sign__12_comb = p2_is_operand_inf__1 ? p2_not_5126 : p3_result_sign__11_comb;
  assign p3_rounded_fraction_comb = p3_do_round_up__5_comb ? {p3_add_5248_comb, p3_normal_chunk_comb} : {1'h0, p3_shifted_fraction_comb};
  assign p3_rounded_fraction__1_comb = p3_do_round_up__6_comb ? {p3_add_5252_comb, p3_normal_chunk__1_comb} : {1'h0, p3_shifted_fraction__1_comb};
  assign p3_ne_5263_comb = p3_fraction__33_comb != 29'h0000_0000;
  assign p3_ne_5264_comb = p3_fraction__34_comb != 29'h0000_0000;
  assign p3_result_sign__13_comb = ~p2_is_result_nan__5 & p3_result_sign__10_comb;
  assign p3_result_sign__14_comb = ~p2_is_result_nan__6 & p3_result_sign__12_comb;

  // Registers for pipe stage 3:
  reg [7:0] p3_greater_exp_bexp;
  reg [7:0] p3_greater_exp_bexp__1;
  reg [4:0] p3_encode_5179;
  reg [4:0] p3_encode_5180;
  reg [27:0] p3_rounded_fraction;
  reg [27:0] p3_rounded_fraction__1;
  reg p3_ne_5263;
  reg p3_ne_5264;
  reg p3_nor_5116;
  reg p3_nor_5120;
  reg p3_is_result_nan__5;
  reg p3_is_operand_inf;
  reg p3_is_result_nan__6;
  reg p3_is_operand_inf__1;
  reg p3_result_sign__13;
  reg p3_result_sign__14;
  always_ff @ (posedge clk) begin
    p3_greater_exp_bexp <= p2_greater_exp_bexp;
    p3_greater_exp_bexp__1 <= p2_greater_exp_bexp__1;
    p3_encode_5179 <= p3_encode_5179_comb;
    p3_encode_5180 <= p3_encode_5180_comb;
    p3_rounded_fraction <= p3_rounded_fraction_comb;
    p3_rounded_fraction__1 <= p3_rounded_fraction__1_comb;
    p3_ne_5263 <= p3_ne_5263_comb;
    p3_ne_5264 <= p3_ne_5264_comb;
    p3_nor_5116 <= p2_nor_5116;
    p3_nor_5120 <= p2_nor_5120;
    p3_is_result_nan__5 <= p2_is_result_nan__5;
    p3_is_operand_inf <= p2_is_operand_inf;
    p3_is_result_nan__6 <= p2_is_result_nan__6;
    p3_is_operand_inf__1 <= p2_is_operand_inf__1;
    p3_result_sign__13 <= p3_result_sign__13_comb;
    p3_result_sign__14 <= p3_result_sign__14_comb;
  end

  // ===== Pipe stage 4:
  wire p4_rounding_carry_comb;
  wire p4_rounding_carry__1_comb;
  wire [8:0] p4_add_5332_comb;
  wire [8:0] p4_add_5334_comb;
  wire [9:0] p4_add_5341_comb;
  wire [9:0] p4_add_5343_comb;
  wire [9:0] p4_wide_exponent_comb;
  wire [9:0] p4_wide_exponent__3_comb;
  wire [9:0] p4_wide_exponent__1_comb;
  wire [9:0] p4_wide_exponent__4_comb;
  wire [8:0] p4_wide_exponent__2_comb;
  wire [8:0] p4_wide_exponent__5_comb;
  wire [2:0] p4_add_5388_comb;
  wire [2:0] p4_add_5391_comb;
  wire p4_nor_5393_comb;
  wire [27:0] p4_shrl_5394_comb;
  wire p4_nor_5396_comb;
  wire [27:0] p4_shrl_5397_comb;
  wire [22:0] p4_result_fraction__13_comb;
  wire [22:0] p4_result_fraction__15_comb;
  wire [7:0] p4_high_exp__26_comb;
  wire [22:0] p4_result_fraction__14_comb;
  wire [22:0] p4_nan_fraction__10_comb;
  wire [7:0] p4_high_exp__27_comb;
  wire [22:0] p4_result_fraction__16_comb;
  wire [22:0] p4_nan_fraction__11_comb;
  wire [7:0] p4_result_exponent__2_comb;
  wire [22:0] p4_result_fraction__17_comb;
  wire [7:0] p4_result_exponent__1_comb;
  wire [22:0] p4_result_fraction__18_comb;
  wire [31:0] p4_re_comb;
  wire [31:0] p4_im_comb;
  wire [31:0] p4_array_5425_comb[2];
  assign p4_rounding_carry_comb = p3_rounded_fraction[27];
  assign p4_rounding_carry__1_comb = p3_rounded_fraction__1[27];
  assign p4_add_5332_comb = {1'h0, p3_greater_exp_bexp} + {8'h00, p4_rounding_carry_comb};
  assign p4_add_5334_comb = {1'h0, p3_greater_exp_bexp__1} + {8'h00, p4_rounding_carry__1_comb};
  assign p4_add_5341_comb = {1'h0, p4_add_5332_comb} + 10'h001;
  assign p4_add_5343_comb = {1'h0, p4_add_5334_comb} + 10'h001;
  assign p4_wide_exponent_comb = p4_add_5341_comb - {5'h00, p3_encode_5179};
  assign p4_wide_exponent__3_comb = p4_add_5343_comb - {5'h00, p3_encode_5180};
  assign p4_wide_exponent__1_comb = p4_wide_exponent_comb & {10{p3_ne_5263}};
  assign p4_wide_exponent__4_comb = p4_wide_exponent__3_comb & {10{p3_ne_5264}};
  assign p4_wide_exponent__2_comb = p4_wide_exponent__1_comb[8:0] & {9{~p4_wide_exponent__1_comb[9]}};
  assign p4_wide_exponent__5_comb = p4_wide_exponent__4_comb[8:0] & {9{~p4_wide_exponent__4_comb[9]}};
  assign p4_add_5388_comb = {2'h0, p4_rounding_carry_comb} + 3'h3;
  assign p4_add_5391_comb = {2'h0, p4_rounding_carry__1_comb} + 3'h3;
  assign p4_nor_5393_comb = ~(p4_wide_exponent__2_comb[8] | p4_wide_exponent__2_comb[0] & p4_wide_exponent__2_comb[1] & p4_wide_exponent__2_comb[2] & p4_wide_exponent__2_comb[3] & p4_wide_exponent__2_comb[4] & p4_wide_exponent__2_comb[5] & p4_wide_exponent__2_comb[6] & p4_wide_exponent__2_comb[7]);
  assign p4_shrl_5394_comb = p3_rounded_fraction >> p4_add_5388_comb;
  assign p4_nor_5396_comb = ~(p4_wide_exponent__5_comb[8] | p4_wide_exponent__5_comb[0] & p4_wide_exponent__5_comb[1] & p4_wide_exponent__5_comb[2] & p4_wide_exponent__5_comb[3] & p4_wide_exponent__5_comb[4] & p4_wide_exponent__5_comb[5] & p4_wide_exponent__5_comb[6] & p4_wide_exponent__5_comb[7]);
  assign p4_shrl_5397_comb = p3_rounded_fraction__1 >> p4_add_5391_comb;
  assign p4_result_fraction__13_comb = p4_shrl_5394_comb[22:0];
  assign p4_result_fraction__15_comb = p4_shrl_5397_comb[22:0];
  assign p4_high_exp__26_comb = 8'hff;
  assign p4_result_fraction__14_comb = p4_result_fraction__13_comb & {23{~(~(p4_wide_exponent__2_comb[1] | p4_wide_exponent__2_comb[2] | p4_wide_exponent__2_comb[3] | p4_wide_exponent__2_comb[4] | p4_wide_exponent__2_comb[5] | p4_wide_exponent__2_comb[6] | p4_wide_exponent__2_comb[7] | p4_wide_exponent__2_comb[8] | p4_wide_exponent__2_comb[0]))}} & {23{p4_nor_5393_comb}} & {23{p3_nor_5116}};
  assign p4_nan_fraction__10_comb = 23'h40_0000;
  assign p4_high_exp__27_comb = 8'hff;
  assign p4_result_fraction__16_comb = p4_result_fraction__15_comb & {23{~(~(p4_wide_exponent__5_comb[1] | p4_wide_exponent__5_comb[2] | p4_wide_exponent__5_comb[3] | p4_wide_exponent__5_comb[4] | p4_wide_exponent__5_comb[5] | p4_wide_exponent__5_comb[6] | p4_wide_exponent__5_comb[7] | p4_wide_exponent__5_comb[8] | p4_wide_exponent__5_comb[0]))}} & {23{p4_nor_5396_comb}} & {23{p3_nor_5120}};
  assign p4_nan_fraction__11_comb = 23'h40_0000;
  assign p4_result_exponent__2_comb = p3_is_result_nan__5 | p3_is_operand_inf | ~p4_nor_5393_comb ? p4_high_exp__26_comb : p4_wide_exponent__2_comb[7:0];
  assign p4_result_fraction__17_comb = p3_is_result_nan__5 ? p4_nan_fraction__10_comb : p4_result_fraction__14_comb;
  assign p4_result_exponent__1_comb = p3_is_result_nan__6 | p3_is_operand_inf__1 | ~p4_nor_5396_comb ? p4_high_exp__27_comb : p4_wide_exponent__5_comb[7:0];
  assign p4_result_fraction__18_comb = p3_is_result_nan__6 ? p4_nan_fraction__11_comb : p4_result_fraction__16_comb;
  assign p4_re_comb = {p3_result_sign__13, p4_result_exponent__2_comb, p4_result_fraction__17_comb};
  assign p4_im_comb = {p3_result_sign__14, p4_result_exponent__1_comb, p4_result_fraction__18_comb};
  assign p4_array_5425_comb[0] = p4_re_comb;
  assign p4_array_5425_comb[1] = p4_im_comb;

  // Registers for pipe stage 4:
  reg [31:0] p4_array_5425[2];
  always_ff @ (posedge clk) begin
    p4_array_5425 <= p4_array_5425_comb;
  end
  __tmp__ComplexMult_17___itok__tmp__ComplexMult___itok__tmp__ComplexMult_15___itok__apfloat__sub__8_23___itok__apfloat__sub__8_23_10___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p3_and_5209_comb | p3_and_5208_comb | p3_and_5207_comb)) p3_and_5209_comb | p3_and_5208_comb | p3_and_5207_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  __tmp__ComplexMult_17___itok__tmp__ComplexMult___itok__tmp__ComplexMult_16___itok__apfloat__add__8_23_carry_and_cancel: assert property (@(posedge clk) disable iff ($isunknown(p3_and_5216_comb | p3_and_5215_comb | p3_and_5214_comb)) p3_and_5216_comb | p3_and_5215_comb | p3_and_5214_comb) else $fatal(0, "Assertion failure via fail! @ xls/dslx/stdlib/apfloat.x:1683:15-1683:62");
  assign out = {p4_array_5425[1], p4_array_5425[0]};
endmodule
